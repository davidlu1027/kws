`timescale 1ns/10ps

module fft_r22sdf_rom_1024_s2 (
    input  wire               clk,
    input  wire               rst_n,
    input  wire        [ 5:0] addr,
    input  wire               addr_vld,
    output reg signed [ 9:0] tf_re,
    output reg signed [ 9:0] tf_im
  );

  reg  [19:0] dout[0:63];

  // assign tf_re = dout[19:10];
  // assign tf_im = dout[ 9: 0];

  // initial
  //   begin
  //    `ifndef USE_RESET
  //     dout = 20'd0;
  //    `endif
  //   end

  // always @ (posedge clk or negedge rst_n)
  //   begin
  //     if (!rst_n)
  //       begin
  //       //  `ifdef USE_RESET
  //         dout <= 20'd0;
  //       //  `endif
  //       end
  //     else if (addr_vld)
  //       begin
  //         case (addr)
initial begin
dout[0]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[1]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[2]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[3]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[4]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[5]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[6]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[7]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[8]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[9]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[10]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[11]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[12]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[13]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[14]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[15]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[16]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[17]=	{ 10'sd502   , -10'sd100   }; /* W[  32] =  0.9805  -0.1953i */
dout[18]=	{ 10'sd473   , -10'sd196   }; /* W[  64] =  0.9238  -0.3828i */
dout[19]=	{ 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[20]=	{ 10'sd362   , -10'sd362   }; /* W[ 128] =  0.7070  -0.7070i */
dout[21]=	{ 10'sd284   , -10'sd426   }; /* W[ 160] =  0.5547  -0.8320i */
dout[22]=	{ 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[23]=	{ 10'sd100   , -10'sd502   }; /* W[ 224] =  0.1953  -0.9805i */
dout[24]=	{ 10'sd0     , -10'sd512   }; /* W[ 256] =  0.0000  -1.0000i */
dout[25]=	{-10'sd100   , -10'sd502   }; /* W[ 288] = -0.1953  -0.9805i */
dout[26]=	{-10'sd196   , -10'sd473   }; /* W[ 320] = -0.3828  -0.9238i */
dout[27]=	{-10'sd284   , -10'sd426   }; /* W[ 352] = -0.5547  -0.8320i */
dout[28]=	{-10'sd362   , -10'sd362   }; /* W[ 384] = -0.7070  -0.7070i */
dout[29]=	{-10'sd426   , -10'sd284   }; /* W[ 416] = -0.8320  -0.5547i */
dout[30]=	{-10'sd473   , -10'sd196   }; /* W[ 448] = -0.9238  -0.3828i */
dout[31]=	{-10'sd502   , -10'sd100   }; /* W[ 480] = -0.9805  -0.1953i */
dout[32]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[33]=	{ 10'sd510   , -10'sd50    }; /* W[  16] =  0.9961  -0.0977i */
dout[34]=	{ 10'sd502   , -10'sd100   }; /* W[  32] =  0.9805  -0.1953i */
dout[35]=	{ 10'sd490   , -10'sd149   }; /* W[  48] =  0.9570  -0.2910i */
dout[36]=	{ 10'sd473   , -10'sd196   }; /* W[  64] =  0.9238  -0.3828i */
dout[37]=	{ 10'sd452   , -10'sd241   }; /* W[  80] =  0.8828  -0.4707i */
dout[38]=	{ 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[39]=	{ 10'sd396   , -10'sd325   }; /* W[ 112] =  0.7734  -0.6348i */
dout[40]=	{ 10'sd362   , -10'sd362   }; /* W[ 128] =  0.7070  -0.7070i */
dout[41]=	{ 10'sd325   , -10'sd396   }; /* W[ 144] =  0.6348  -0.7734i */
dout[42]=	{ 10'sd284   , -10'sd426   }; /* W[ 160] =  0.5547  -0.8320i */
dout[43]=	{ 10'sd241   , -10'sd452   }; /* W[ 176] =  0.4707  -0.8828i */
dout[44]=	{ 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[45]=	{ 10'sd149   , -10'sd490   }; /* W[ 208] =  0.2910  -0.9570i */
dout[46]=	{ 10'sd100   , -10'sd502   }; /* W[ 224] =  0.1953  -0.9805i */
dout[47]=	{ 10'sd50    , -10'sd510   }; /* W[ 240] =  0.0977  -0.9961i */
dout[48]=	{ 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[49]=	{ 10'sd490   , -10'sd149   }; /* W[  48] =  0.9570  -0.2910i */
dout[50]=	{ 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[51]=	{ 10'sd325   , -10'sd396   }; /* W[ 144] =  0.6348  -0.7734i */
dout[52]=	{ 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[53]=	{ 10'sd50    , -10'sd510   }; /* W[ 240] =  0.0977  -0.9961i */
dout[54]=	{-10'sd100   , -10'sd502   }; /* W[ 288] = -0.1953  -0.9805i */
dout[55]=	{-10'sd241   , -10'sd452   }; /* W[ 336] = -0.4707  -0.8828i */
dout[56]=	{-10'sd362   , -10'sd362   }; /* W[ 384] = -0.7070  -0.7070i */
dout[57]=	{-10'sd452   , -10'sd241   }; /* W[ 432] = -0.8828  -0.4707i */
dout[58]=	{-10'sd502   , -10'sd100   }; /* W[ 480] = -0.9805  -0.1953i */
dout[59]=	{-10'sd510   ,  10'sd50    }; /* W[ 528] = -0.9961   0.0977i */
dout[60]=	{-10'sd473   ,  10'sd196   }; /* W[ 576] = -0.9238   0.3828i */
dout[61]=	{-10'sd396   ,  10'sd325   }; /* W[ 624] = -0.7734   0.6348i */
dout[62]=	{-10'sd284   ,  10'sd426   }; /* W[ 672] = -0.5547   0.8320i */
dout[63]=	{-10'sd149   ,  10'sd490   }; /* W[ 720] = -0.2910   0.9570i */
end

always @ (posedge clk) begin
  tf_re<=dout[addr][19:10];
  tf_im<=dout[addr][9:0];
end


endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */
