module hamming_window_rom (
    input  wire               clk,
    input  wire               rst_n,
    input  wire        [ 9:0] addr,
    input  wire               in_valid,
    output reg signed [ 11:0] w
  );
reg  [11:0] dout[0:1023];

initial begin
dout[0]=12'd327;
dout[1]=12'd327;
dout[2]=12'd327;
dout[3]=12'd327;
dout[4]=12'd328;
dout[5]=12'd328;
dout[6]=12'd328;
dout[7]=12'd329;
dout[8]=12'd329;
dout[9]=12'd330;
dout[10]=12'd331;
dout[11]=12'd331;
dout[12]=12'd332;
dout[13]=12'd333;
dout[14]=12'd334;
dout[15]=12'd335;
dout[16]=12'd336;
dout[17]=12'd337;
dout[18]=12'd339;
dout[19]=12'd340;
dout[20]=12'd341;
dout[21]=12'd343;
dout[22]=12'd344;
dout[23]=12'd346;
dout[24]=12'd348;
dout[25]=12'd349;
dout[26]=12'd351;
dout[27]=12'd353;
dout[28]=12'd355;
dout[29]=12'd357;
dout[30]=12'd359;
dout[31]=12'd361;
dout[32]=12'd363;
dout[33]=12'd366;
dout[34]=12'd368;
dout[35]=12'd371;
dout[36]=12'd373;
dout[37]=12'd376;
dout[38]=12'd378;
dout[39]=12'd381;
dout[40]=12'd384;
dout[41]=12'd387;
dout[42]=12'd390;
dout[43]=12'd393;
dout[44]=12'd396;
dout[45]=12'd399;
dout[46]=12'd402;
dout[47]=12'd405;
dout[48]=12'd408;
dout[49]=12'd412;
dout[50]=12'd415;
dout[51]=12'd419;
dout[52]=12'd422;
dout[53]=12'd426;
dout[54]=12'd430;
dout[55]=12'd434;
dout[56]=12'd438;
dout[57]=12'd441;
dout[58]=12'd445;
dout[59]=12'd450;
dout[60]=12'd454;
dout[61]=12'd458;
dout[62]=12'd462;
dout[63]=12'd466;
dout[64]=12'd471;
dout[65]=12'd475;
dout[66]=12'd480;
dout[67]=12'd484;
dout[68]=12'd489;
dout[69]=12'd494;
dout[70]=12'd499;
dout[71]=12'd504;
dout[72]=12'd508;
dout[73]=12'd513;
dout[74]=12'd518;
dout[75]=12'd524;
dout[76]=12'd529;
dout[77]=12'd534;
dout[78]=12'd539;
dout[79]=12'd545;
dout[80]=12'd550;
dout[81]=12'd556;
dout[82]=12'd561;
dout[83]=12'd567;
dout[84]=12'd572;
dout[85]=12'd578;
dout[86]=12'd584;
dout[87]=12'd590;
dout[88]=12'd596;
dout[89]=12'd602;
dout[90]=12'd608;
dout[91]=12'd614;
dout[92]=12'd620;
dout[93]=12'd626;
dout[94]=12'd633;
dout[95]=12'd639;
dout[96]=12'd645;
dout[97]=12'd652;
dout[98]=12'd658;
dout[99]=12'd665;
dout[100]=12'd672;
dout[101]=12'd678;
dout[102]=12'd685;
dout[103]=12'd692;
dout[104]=12'd699;
dout[105]=12'd706;
dout[106]=12'd713;
dout[107]=12'd720;
dout[108]=12'd727;
dout[109]=12'd734;
dout[110]=12'd741;
dout[111]=12'd748;
dout[112]=12'd756;
dout[113]=12'd763;
dout[114]=12'd770;
dout[115]=12'd778;
dout[116]=12'd785;
dout[117]=12'd793;
dout[118]=12'd801;
dout[119]=12'd808;
dout[120]=12'd816;
dout[121]=12'd824;
dout[122]=12'd832;
dout[123]=12'd840;
dout[124]=12'd848;
dout[125]=12'd856;
dout[126]=12'd864;
dout[127]=12'd872;
dout[128]=12'd880;
dout[129]=12'd888;
dout[130]=12'd897;
dout[131]=12'd905;
dout[132]=12'd913;
dout[133]=12'd922;
dout[134]=12'd930;
dout[135]=12'd939;
dout[136]=12'd947;
dout[137]=12'd956;
dout[138]=12'd964;
dout[139]=12'd973;
dout[140]=12'd982;
dout[141]=12'd991;
dout[142]=12'd999;
dout[143]=12'd1008;
dout[144]=12'd1017;
dout[145]=12'd1026;
dout[146]=12'd1035;
dout[147]=12'd1044;
dout[148]=12'd1053;
dout[149]=12'd1063;
dout[150]=12'd1072;
dout[151]=12'd1081;
dout[152]=12'd1090;
dout[153]=12'd1100;
dout[154]=12'd1109;
dout[155]=12'd1118;
dout[156]=12'd1128;
dout[157]=12'd1137;
dout[158]=12'd1147;
dout[159]=12'd1156;
dout[160]=12'd1166;
dout[161]=12'd1176;
dout[162]=12'd1185;
dout[163]=12'd1195;
dout[164]=12'd1205;
dout[165]=12'd1215;
dout[166]=12'd1225;
dout[167]=12'd1234;
dout[168]=12'd1244;
dout[169]=12'd1254;
dout[170]=12'd1264;
dout[171]=12'd1274;
dout[172]=12'd1284;
dout[173]=12'd1294;
dout[174]=12'd1305;
dout[175]=12'd1315;
dout[176]=12'd1325;
dout[177]=12'd1335;
dout[178]=12'd1345;
dout[179]=12'd1356;
dout[180]=12'd1366;
dout[181]=12'd1376;
dout[182]=12'd1387;
dout[183]=12'd1397;
dout[184]=12'd1408;
dout[185]=12'd1418;
dout[186]=12'd1429;
dout[187]=12'd1439;
dout[188]=12'd1450;
dout[189]=12'd1460;
dout[190]=12'd1471;
dout[191]=12'd1482;
dout[192]=12'd1492;
dout[193]=12'd1503;
dout[194]=12'd1514;
dout[195]=12'd1525;
dout[196]=12'd1535;
dout[197]=12'd1546;
dout[198]=12'd1557;
dout[199]=12'd1568;
dout[200]=12'd1579;
dout[201]=12'd1590;
dout[202]=12'd1601;
dout[203]=12'd1612;
dout[204]=12'd1623;
dout[205]=12'd1634;
dout[206]=12'd1645;
dout[207]=12'd1656;
dout[208]=12'd1667;
dout[209]=12'd1678;
dout[210]=12'd1689;
dout[211]=12'd1700;
dout[212]=12'd1711;
dout[213]=12'd1722;
dout[214]=12'd1733;
dout[215]=12'd1745;
dout[216]=12'd1756;
dout[217]=12'd1767;
dout[218]=12'd1778;
dout[219]=12'd1790;
dout[220]=12'd1801;
dout[221]=12'd1812;
dout[222]=12'd1824;
dout[223]=12'd1835;
dout[224]=12'd1846;
dout[225]=12'd1858;
dout[226]=12'd1869;
dout[227]=12'd1880;
dout[228]=12'd1892;
dout[229]=12'd1903;
dout[230]=12'd1915;
dout[231]=12'd1926;
dout[232]=12'd1937;
dout[233]=12'd1949;
dout[234]=12'd1960;
dout[235]=12'd1972;
dout[236]=12'd1983;
dout[237]=12'd1995;
dout[238]=12'd2006;
dout[239]=12'd2018;
dout[240]=12'd2029;
dout[241]=12'd2041;
dout[242]=12'd2052;
dout[243]=12'd2064;
dout[244]=12'd2075;
dout[245]=12'd2087;
dout[246]=12'd2099;
dout[247]=12'd2110;
dout[248]=12'd2122;
dout[249]=12'd2133;
dout[250]=12'd2145;
dout[251]=12'd2156;
dout[252]=12'd2168;
dout[253]=12'd2180;
dout[254]=12'd2191;
dout[255]=12'd2203;
dout[256]=12'd2214;
dout[257]=12'd2226;
dout[258]=12'd2237;
dout[259]=12'd2249;
dout[260]=12'd2261;
dout[261]=12'd2272;
dout[262]=12'd2284;
dout[263]=12'd2295;
dout[264]=12'd2307;
dout[265]=12'd2318;
dout[266]=12'd2330;
dout[267]=12'd2341;
dout[268]=12'd2353;
dout[269]=12'd2365;
dout[270]=12'd2376;
dout[271]=12'd2388;
dout[272]=12'd2399;
dout[273]=12'd2411;
dout[274]=12'd2422;
dout[275]=12'd2434;
dout[276]=12'd2445;
dout[277]=12'd2457;
dout[278]=12'd2468;
dout[279]=12'd2479;
dout[280]=12'd2491;
dout[281]=12'd2502;
dout[282]=12'd2514;
dout[283]=12'd2525;
dout[284]=12'd2537;
dout[285]=12'd2548;
dout[286]=12'd2559;
dout[287]=12'd2571;
dout[288]=12'd2582;
dout[289]=12'd2593;
dout[290]=12'd2605;
dout[291]=12'd2616;
dout[292]=12'd2627;
dout[293]=12'd2639;
dout[294]=12'd2650;
dout[295]=12'd2661;
dout[296]=12'd2672;
dout[297]=12'd2684;
dout[298]=12'd2695;
dout[299]=12'd2706;
dout[300]=12'd2717;
dout[301]=12'd2728;
dout[302]=12'd2739;
dout[303]=12'd2750;
dout[304]=12'd2762;
dout[305]=12'd2773;
dout[306]=12'd2784;
dout[307]=12'd2795;
dout[308]=12'd2806;
dout[309]=12'd2817;
dout[310]=12'd2828;
dout[311]=12'd2839;
dout[312]=12'd2849;
dout[313]=12'd2860;
dout[314]=12'd2871;
dout[315]=12'd2882;
dout[316]=12'd2893;
dout[317]=12'd2904;
dout[318]=12'd2914;
dout[319]=12'd2925;
dout[320]=12'd2936;
dout[321]=12'd2946;
dout[322]=12'd2957;
dout[323]=12'd2968;
dout[324]=12'd2978;
dout[325]=12'd2989;
dout[326]=12'd2999;
dout[327]=12'd3010;
dout[328]=12'd3020;
dout[329]=12'd3031;
dout[330]=12'd3041;
dout[331]=12'd3051;
dout[332]=12'd3062;
dout[333]=12'd3072;
dout[334]=12'd3082;
dout[335]=12'd3093;
dout[336]=12'd3103;
dout[337]=12'd3113;
dout[338]=12'd3123;
dout[339]=12'd3133;
dout[340]=12'd3143;
dout[341]=12'd3153;
dout[342]=12'd3163;
dout[343]=12'd3173;
dout[344]=12'd3183;
dout[345]=12'd3193;
dout[346]=12'd3203;
dout[347]=12'd3213;
dout[348]=12'd3223;
dout[349]=12'd3232;
dout[350]=12'd3242;
dout[351]=12'd3252;
dout[352]=12'd3261;
dout[353]=12'd3271;
dout[354]=12'd3281;
dout[355]=12'd3290;
dout[356]=12'd3300;
dout[357]=12'd3309;
dout[358]=12'd3318;
dout[359]=12'd3328;
dout[360]=12'd3337;
dout[361]=12'd3346;
dout[362]=12'd3355;
dout[363]=12'd3365;
dout[364]=12'd3374;
dout[365]=12'd3383;
dout[366]=12'd3392;
dout[367]=12'd3401;
dout[368]=12'd3410;
dout[369]=12'd3419;
dout[370]=12'd3428;
dout[371]=12'd3436;
dout[372]=12'd3445;
dout[373]=12'd3454;
dout[374]=12'd3463;
dout[375]=12'd3471;
dout[376]=12'd3480;
dout[377]=12'd3488;
dout[378]=12'd3497;
dout[379]=12'd3505;
dout[380]=12'd3514;
dout[381]=12'd3522;
dout[382]=12'd3530;
dout[383]=12'd3539;
dout[384]=12'd3547;
dout[385]=12'd3555;
dout[386]=12'd3563;
dout[387]=12'd3571;
dout[388]=12'd3579;
dout[389]=12'd3587;
dout[390]=12'd3595;
dout[391]=12'd3603;
dout[392]=12'd3610;
dout[393]=12'd3618;
dout[394]=12'd3626;
dout[395]=12'd3633;
dout[396]=12'd3641;
dout[397]=12'd3648;
dout[398]=12'd3656;
dout[399]=12'd3663;
dout[400]=12'd3671;
dout[401]=12'd3678;
dout[402]=12'd3685;
dout[403]=12'd3692;
dout[404]=12'd3700;
dout[405]=12'd3707;
dout[406]=12'd3714;
dout[407]=12'd3721;
dout[408]=12'd3727;
dout[409]=12'd3734;
dout[410]=12'd3741;
dout[411]=12'd3748;
dout[412]=12'd3754;
dout[413]=12'd3761;
dout[414]=12'd3768;
dout[415]=12'd3774;
dout[416]=12'd3781;
dout[417]=12'd3787;
dout[418]=12'd3793;
dout[419]=12'd3800;
dout[420]=12'd3806;
dout[421]=12'd3812;
dout[422]=12'd3818;
dout[423]=12'd3824;
dout[424]=12'd3830;
dout[425]=12'd3836;
dout[426]=12'd3842;
dout[427]=12'd3847;
dout[428]=12'd3853;
dout[429]=12'd3859;
dout[430]=12'd3864;
dout[431]=12'd3870;
dout[432]=12'd3875;
dout[433]=12'd3881;
dout[434]=12'd3886;
dout[435]=12'd3891;
dout[436]=12'd3897;
dout[437]=12'd3902;
dout[438]=12'd3907;
dout[439]=12'd3912;
dout[440]=12'd3917;
dout[441]=12'd3922;
dout[442]=12'd3926;
dout[443]=12'd3931;
dout[444]=12'd3936;
dout[445]=12'd3941;
dout[446]=12'd3945;
dout[447]=12'd3950;
dout[448]=12'd3954;
dout[449]=12'd3958;
dout[450]=12'd3963;
dout[451]=12'd3967;
dout[452]=12'd3971;
dout[453]=12'd3975;
dout[454]=12'd3979;
dout[455]=12'd3983;
dout[456]=12'd3987;
dout[457]=12'd3991;
dout[458]=12'd3995;
dout[459]=12'd3998;
dout[460]=12'd4002;
dout[461]=12'd4006;
dout[462]=12'd4009;
dout[463]=12'd4013;
dout[464]=12'd4016;
dout[465]=12'd4019;
dout[466]=12'd4022;
dout[467]=12'd4026;
dout[468]=12'd4029;
dout[469]=12'd4032;
dout[470]=12'd4035;
dout[471]=12'd4038;
dout[472]=12'd4040;
dout[473]=12'd4043;
dout[474]=12'd4046;
dout[475]=12'd4048;
dout[476]=12'd4051;
dout[477]=12'd4053;
dout[478]=12'd4056;
dout[479]=12'd4058;
dout[480]=12'd4060;
dout[481]=12'd4063;
dout[482]=12'd4065;
dout[483]=12'd4067;
dout[484]=12'd4069;
dout[485]=12'd4071;
dout[486]=12'd4072;
dout[487]=12'd4074;
dout[488]=12'd4076;
dout[489]=12'd4078;
dout[490]=12'd4079;
dout[491]=12'd4081;
dout[492]=12'd4082;
dout[493]=12'd4083;
dout[494]=12'd4085;
dout[495]=12'd4086;
dout[496]=12'd4087;
dout[497]=12'd4088;
dout[498]=12'd4089;
dout[499]=12'd4090;
dout[500]=12'd4091;
dout[501]=12'd4092;
dout[502]=12'd4092;
dout[503]=12'd4093;
dout[504]=12'd4094;
dout[505]=12'd4094;
dout[506]=12'd4094;
dout[507]=12'd4095;
dout[508]=12'd4095;
dout[509]=12'd4095;
dout[510]=12'd4095;
dout[511]=12'd4095;
dout[512]=12'd4095;
dout[513]=12'd4095;
dout[514]=12'd4095;
dout[515]=12'd4095;
dout[516]=12'd4095;
dout[517]=12'd4094;
dout[518]=12'd4094;
dout[519]=12'd4094;
dout[520]=12'd4093;
dout[521]=12'd4092;
dout[522]=12'd4092;
dout[523]=12'd4091;
dout[524]=12'd4090;
dout[525]=12'd4089;
dout[526]=12'd4088;
dout[527]=12'd4087;
dout[528]=12'd4086;
dout[529]=12'd4085;
dout[530]=12'd4083;
dout[531]=12'd4082;
dout[532]=12'd4081;
dout[533]=12'd4079;
dout[534]=12'd4078;
dout[535]=12'd4076;
dout[536]=12'd4074;
dout[537]=12'd4072;
dout[538]=12'd4071;
dout[539]=12'd4069;
dout[540]=12'd4067;
dout[541]=12'd4065;
dout[542]=12'd4063;
dout[543]=12'd4060;
dout[544]=12'd4058;
dout[545]=12'd4056;
dout[546]=12'd4053;
dout[547]=12'd4051;
dout[548]=12'd4048;
dout[549]=12'd4046;
dout[550]=12'd4043;
dout[551]=12'd4040;
dout[552]=12'd4038;
dout[553]=12'd4035;
dout[554]=12'd4032;
dout[555]=12'd4029;
dout[556]=12'd4026;
dout[557]=12'd4022;
dout[558]=12'd4019;
dout[559]=12'd4016;
dout[560]=12'd4013;
dout[561]=12'd4009;
dout[562]=12'd4006;
dout[563]=12'd4002;
dout[564]=12'd3998;
dout[565]=12'd3995;
dout[566]=12'd3991;
dout[567]=12'd3987;
dout[568]=12'd3983;
dout[569]=12'd3979;
dout[570]=12'd3975;
dout[571]=12'd3971;
dout[572]=12'd3967;
dout[573]=12'd3963;
dout[574]=12'd3958;
dout[575]=12'd3954;
dout[576]=12'd3950;
dout[577]=12'd3945;
dout[578]=12'd3941;
dout[579]=12'd3936;
dout[580]=12'd3931;
dout[581]=12'd3926;
dout[582]=12'd3922;
dout[583]=12'd3917;
dout[584]=12'd3912;
dout[585]=12'd3907;
dout[586]=12'd3902;
dout[587]=12'd3897;
dout[588]=12'd3891;
dout[589]=12'd3886;
dout[590]=12'd3881;
dout[591]=12'd3875;
dout[592]=12'd3870;
dout[593]=12'd3864;
dout[594]=12'd3859;
dout[595]=12'd3853;
dout[596]=12'd3847;
dout[597]=12'd3842;
dout[598]=12'd3836;
dout[599]=12'd3830;
dout[600]=12'd3824;
dout[601]=12'd3818;
dout[602]=12'd3812;
dout[603]=12'd3806;
dout[604]=12'd3800;
dout[605]=12'd3793;
dout[606]=12'd3787;
dout[607]=12'd3781;
dout[608]=12'd3774;
dout[609]=12'd3768;
dout[610]=12'd3761;
dout[611]=12'd3754;
dout[612]=12'd3748;
dout[613]=12'd3741;
dout[614]=12'd3734;
dout[615]=12'd3727;
dout[616]=12'd3721;
dout[617]=12'd3714;
dout[618]=12'd3707;
dout[619]=12'd3700;
dout[620]=12'd3692;
dout[621]=12'd3685;
dout[622]=12'd3678;
dout[623]=12'd3671;
dout[624]=12'd3663;
dout[625]=12'd3656;
dout[626]=12'd3648;
dout[627]=12'd3641;
dout[628]=12'd3633;
dout[629]=12'd3626;
dout[630]=12'd3618;
dout[631]=12'd3610;
dout[632]=12'd3603;
dout[633]=12'd3595;
dout[634]=12'd3587;
dout[635]=12'd3579;
dout[636]=12'd3571;
dout[637]=12'd3563;
dout[638]=12'd3555;
dout[639]=12'd3547;
dout[640]=12'd3539;
dout[641]=12'd3530;
dout[642]=12'd3522;
dout[643]=12'd3514;
dout[644]=12'd3505;
dout[645]=12'd3497;
dout[646]=12'd3488;
dout[647]=12'd3480;
dout[648]=12'd3471;
dout[649]=12'd3463;
dout[650]=12'd3454;
dout[651]=12'd3445;
dout[652]=12'd3436;
dout[653]=12'd3428;
dout[654]=12'd3419;
dout[655]=12'd3410;
dout[656]=12'd3401;
dout[657]=12'd3392;
dout[658]=12'd3383;
dout[659]=12'd3374;
dout[660]=12'd3365;
dout[661]=12'd3355;
dout[662]=12'd3346;
dout[663]=12'd3337;
dout[664]=12'd3328;
dout[665]=12'd3318;
dout[666]=12'd3309;
dout[667]=12'd3300;
dout[668]=12'd3290;
dout[669]=12'd3281;
dout[670]=12'd3271;
dout[671]=12'd3261;
dout[672]=12'd3252;
dout[673]=12'd3242;
dout[674]=12'd3232;
dout[675]=12'd3223;
dout[676]=12'd3213;
dout[677]=12'd3203;
dout[678]=12'd3193;
dout[679]=12'd3183;
dout[680]=12'd3173;
dout[681]=12'd3163;
dout[682]=12'd3153;
dout[683]=12'd3143;
dout[684]=12'd3133;
dout[685]=12'd3123;
dout[686]=12'd3113;
dout[687]=12'd3103;
dout[688]=12'd3093;
dout[689]=12'd3082;
dout[690]=12'd3072;
dout[691]=12'd3062;
dout[692]=12'd3051;
dout[693]=12'd3041;
dout[694]=12'd3031;
dout[695]=12'd3020;
dout[696]=12'd3010;
dout[697]=12'd2999;
dout[698]=12'd2989;
dout[699]=12'd2978;
dout[700]=12'd2968;
dout[701]=12'd2957;
dout[702]=12'd2946;
dout[703]=12'd2936;
dout[704]=12'd2925;
dout[705]=12'd2914;
dout[706]=12'd2904;
dout[707]=12'd2893;
dout[708]=12'd2882;
dout[709]=12'd2871;
dout[710]=12'd2860;
dout[711]=12'd2849;
dout[712]=12'd2839;
dout[713]=12'd2828;
dout[714]=12'd2817;
dout[715]=12'd2806;
dout[716]=12'd2795;
dout[717]=12'd2784;
dout[718]=12'd2773;
dout[719]=12'd2762;
dout[720]=12'd2750;
dout[721]=12'd2739;
dout[722]=12'd2728;
dout[723]=12'd2717;
dout[724]=12'd2706;
dout[725]=12'd2695;
dout[726]=12'd2684;
dout[727]=12'd2672;
dout[728]=12'd2661;
dout[729]=12'd2650;
dout[730]=12'd2639;
dout[731]=12'd2627;
dout[732]=12'd2616;
dout[733]=12'd2605;
dout[734]=12'd2593;
dout[735]=12'd2582;
dout[736]=12'd2571;
dout[737]=12'd2559;
dout[738]=12'd2548;
dout[739]=12'd2537;
dout[740]=12'd2525;
dout[741]=12'd2514;
dout[742]=12'd2502;
dout[743]=12'd2491;
dout[744]=12'd2479;
dout[745]=12'd2468;
dout[746]=12'd2457;
dout[747]=12'd2445;
dout[748]=12'd2434;
dout[749]=12'd2422;
dout[750]=12'd2411;
dout[751]=12'd2399;
dout[752]=12'd2388;
dout[753]=12'd2376;
dout[754]=12'd2365;
dout[755]=12'd2353;
dout[756]=12'd2341;
dout[757]=12'd2330;
dout[758]=12'd2318;
dout[759]=12'd2307;
dout[760]=12'd2295;
dout[761]=12'd2284;
dout[762]=12'd2272;
dout[763]=12'd2261;
dout[764]=12'd2249;
dout[765]=12'd2237;
dout[766]=12'd2226;
dout[767]=12'd2214;
dout[768]=12'd2203;
dout[769]=12'd2191;
dout[770]=12'd2180;
dout[771]=12'd2168;
dout[772]=12'd2156;
dout[773]=12'd2145;
dout[774]=12'd2133;
dout[775]=12'd2122;
dout[776]=12'd2110;
dout[777]=12'd2099;
dout[778]=12'd2087;
dout[779]=12'd2075;
dout[780]=12'd2064;
dout[781]=12'd2052;
dout[782]=12'd2041;
dout[783]=12'd2029;
dout[784]=12'd2018;
dout[785]=12'd2006;
dout[786]=12'd1995;
dout[787]=12'd1983;
dout[788]=12'd1972;
dout[789]=12'd1960;
dout[790]=12'd1949;
dout[791]=12'd1937;
dout[792]=12'd1926;
dout[793]=12'd1915;
dout[794]=12'd1903;
dout[795]=12'd1892;
dout[796]=12'd1880;
dout[797]=12'd1869;
dout[798]=12'd1858;
dout[799]=12'd1846;
dout[800]=12'd1835;
dout[801]=12'd1824;
dout[802]=12'd1812;
dout[803]=12'd1801;
dout[804]=12'd1790;
dout[805]=12'd1778;
dout[806]=12'd1767;
dout[807]=12'd1756;
dout[808]=12'd1745;
dout[809]=12'd1733;
dout[810]=12'd1722;
dout[811]=12'd1711;
dout[812]=12'd1700;
dout[813]=12'd1689;
dout[814]=12'd1678;
dout[815]=12'd1667;
dout[816]=12'd1656;
dout[817]=12'd1645;
dout[818]=12'd1634;
dout[819]=12'd1623;
dout[820]=12'd1612;
dout[821]=12'd1601;
dout[822]=12'd1590;
dout[823]=12'd1579;
dout[824]=12'd1568;
dout[825]=12'd1557;
dout[826]=12'd1546;
dout[827]=12'd1535;
dout[828]=12'd1525;
dout[829]=12'd1514;
dout[830]=12'd1503;
dout[831]=12'd1492;
dout[832]=12'd1482;
dout[833]=12'd1471;
dout[834]=12'd1460;
dout[835]=12'd1450;
dout[836]=12'd1439;
dout[837]=12'd1429;
dout[838]=12'd1418;
dout[839]=12'd1408;
dout[840]=12'd1397;
dout[841]=12'd1387;
dout[842]=12'd1376;
dout[843]=12'd1366;
dout[844]=12'd1356;
dout[845]=12'd1345;
dout[846]=12'd1335;
dout[847]=12'd1325;
dout[848]=12'd1315;
dout[849]=12'd1305;
dout[850]=12'd1294;
dout[851]=12'd1284;
dout[852]=12'd1274;
dout[853]=12'd1264;
dout[854]=12'd1254;
dout[855]=12'd1244;
dout[856]=12'd1234;
dout[857]=12'd1225;
dout[858]=12'd1215;
dout[859]=12'd1205;
dout[860]=12'd1195;
dout[861]=12'd1185;
dout[862]=12'd1176;
dout[863]=12'd1166;
dout[864]=12'd1156;
dout[865]=12'd1147;
dout[866]=12'd1137;
dout[867]=12'd1128;
dout[868]=12'd1118;
dout[869]=12'd1109;
dout[870]=12'd1100;
dout[871]=12'd1090;
dout[872]=12'd1081;
dout[873]=12'd1072;
dout[874]=12'd1063;
dout[875]=12'd1053;
dout[876]=12'd1044;
dout[877]=12'd1035;
dout[878]=12'd1026;
dout[879]=12'd1017;
dout[880]=12'd1008;
dout[881]=12'd999;
dout[882]=12'd991;
dout[883]=12'd982;
dout[884]=12'd973;
dout[885]=12'd964;
dout[886]=12'd956;
dout[887]=12'd947;
dout[888]=12'd939;
dout[889]=12'd930;
dout[890]=12'd922;
dout[891]=12'd913;
dout[892]=12'd905;
dout[893]=12'd897;
dout[894]=12'd888;
dout[895]=12'd880;
dout[896]=12'd872;
dout[897]=12'd864;
dout[898]=12'd856;
dout[899]=12'd848;
dout[900]=12'd840;
dout[901]=12'd832;
dout[902]=12'd824;
dout[903]=12'd816;
dout[904]=12'd808;
dout[905]=12'd801;
dout[906]=12'd793;
dout[907]=12'd785;
dout[908]=12'd778;
dout[909]=12'd770;
dout[910]=12'd763;
dout[911]=12'd756;
dout[912]=12'd748;
dout[913]=12'd741;
dout[914]=12'd734;
dout[915]=12'd727;
dout[916]=12'd720;
dout[917]=12'd713;
dout[918]=12'd706;
dout[919]=12'd699;
dout[920]=12'd692;
dout[921]=12'd685;
dout[922]=12'd678;
dout[923]=12'd672;
dout[924]=12'd665;
dout[925]=12'd658;
dout[926]=12'd652;
dout[927]=12'd645;
dout[928]=12'd639;
dout[929]=12'd633;
dout[930]=12'd626;
dout[931]=12'd620;
dout[932]=12'd614;
dout[933]=12'd608;
dout[934]=12'd602;
dout[935]=12'd596;
dout[936]=12'd590;
dout[937]=12'd584;
dout[938]=12'd578;
dout[939]=12'd572;
dout[940]=12'd567;
dout[941]=12'd561;
dout[942]=12'd556;
dout[943]=12'd550;
dout[944]=12'd545;
dout[945]=12'd539;
dout[946]=12'd534;
dout[947]=12'd529;
dout[948]=12'd524;
dout[949]=12'd518;
dout[950]=12'd513;
dout[951]=12'd508;
dout[952]=12'd504;
dout[953]=12'd499;
dout[954]=12'd494;
dout[955]=12'd489;
dout[956]=12'd484;
dout[957]=12'd480;
dout[958]=12'd475;
dout[959]=12'd471;
dout[960]=12'd466;
dout[961]=12'd462;
dout[962]=12'd458;
dout[963]=12'd454;
dout[964]=12'd450;
dout[965]=12'd445;
dout[966]=12'd441;
dout[967]=12'd438;
dout[968]=12'd434;
dout[969]=12'd430;
dout[970]=12'd426;
dout[971]=12'd422;
dout[972]=12'd419;
dout[973]=12'd415;
dout[974]=12'd412;
dout[975]=12'd408;
dout[976]=12'd405;
dout[977]=12'd402;
dout[978]=12'd399;
dout[979]=12'd396;
dout[980]=12'd393;
dout[981]=12'd390;
dout[982]=12'd387;
dout[983]=12'd384;
dout[984]=12'd381;
dout[985]=12'd378;
dout[986]=12'd376;
dout[987]=12'd373;
dout[988]=12'd371;
dout[989]=12'd368;
dout[990]=12'd366;
dout[991]=12'd363;
dout[992]=12'd361;
dout[993]=12'd359;
dout[994]=12'd357;
dout[995]=12'd355;
dout[996]=12'd353;
dout[997]=12'd351;
dout[998]=12'd349;
dout[999]=12'd348;
dout[1000]=12'd346;
dout[1001]=12'd344;
dout[1002]=12'd343;
dout[1003]=12'd341;
dout[1004]=12'd340;
dout[1005]=12'd339;
dout[1006]=12'd337;
dout[1007]=12'd336;
dout[1008]=12'd335;
dout[1009]=12'd334;
dout[1010]=12'd333;
dout[1011]=12'd332;
dout[1012]=12'd331;
dout[1013]=12'd331;
dout[1014]=12'd330;
dout[1015]=12'd329;
dout[1016]=12'd329;
dout[1017]=12'd328;
dout[1018]=12'd328;
dout[1019]=12'd328;
dout[1020]=12'd327;
dout[1021]=12'd327;
dout[1022]=12'd327;
dout[1023]=12'd327;
end
always @ (posedge clk) begin
  w <= dout[addr];
end


endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */
