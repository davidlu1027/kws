`timescale 1ns/10ps
module fft_r22sdf_rom_1024_s0 (
    input  wire               clk,
    input  wire               rst_n,
    input  wire        [ 9:0] addr,
    input  wire               addr_vld,
    output reg signed [ 9:0] tf_re,
    output reg signed [ 9:0] tf_im
  );

  reg  [19:0] dout[0:1023];


initial begin
dout[0]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[1]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[2]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[3]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[4]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[5]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[6]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[7]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[8]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[9]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[10]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[11]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[12]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[13]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[14]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[15]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[16]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[17]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[18]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[19]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[20]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[21]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[22]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[23]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[24]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[25]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[26]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[27]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[28]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[29]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[30]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[31]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[32]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[33]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[34]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[35]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[36]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[37]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[38]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[39]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[40]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[41]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[42]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[43]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[44]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[45]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[46]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[47]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[48]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[49]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[50]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[51]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[52]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[53]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[54]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[55]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[56]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[57]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[58]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[59]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[60]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[61]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[62]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[63]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[64]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[65]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[66]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[67]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[68]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[69]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[70]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[71]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[72]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[73]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[74]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[75]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[76]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[77]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[78]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[79]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[80]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[81]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[82]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[83]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[84]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[85]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[86]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[87]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[88]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[89]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[90]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[91]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[92]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[93]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[94]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[95]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[96]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[97]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[98]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[99]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[100]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[101]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[102]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[103]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[104]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[105]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[106]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[107]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[108]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[109]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[110]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[111]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[112]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[113]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[114]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[115]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[116]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[117]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[118]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[119]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[120]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[121]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[122]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[123]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[124]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[125]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[126]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[127]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[128]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[129]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[130]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[131]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[132]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[133]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[134]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[135]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[136]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[137]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[138]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[139]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[140]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[141]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[142]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[143]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[144]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[145]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[146]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[147]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[148]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[149]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[150]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[151]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[152]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[153]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[154]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[155]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[156]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[157]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[158]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[159]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[160]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[161]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[162]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[163]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[164]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[165]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[166]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[167]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[168]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[169]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[170]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[171]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[172]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[173]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[174]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[175]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[176]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[177]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[178]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[179]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[180]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[181]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[182]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[183]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[184]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[185]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[186]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[187]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[188]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[189]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[190]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[191]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[192]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[193]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[194]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[195]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[196]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[197]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[198]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[199]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[200]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[201]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[202]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[203]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[204]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[205]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[206]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[207]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[208]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[209]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[210]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[211]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[212]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[213]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[214]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[215]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[216]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[217]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[218]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[219]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[220]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[221]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[222]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[223]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[224]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[225]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[226]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[227]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[228]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[229]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[230]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[231]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[232]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[233]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[234]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[235]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[236]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[237]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[238]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[239]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[240]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[241]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[242]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[243]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[244]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[245]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[246]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[247]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[248]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[249]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[250]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[251]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[252]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[253]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[254]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[255]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[256]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[257]= { 10'sd511   , -10'sd6     }; /* W[   2] =  0.9980  -0.0117i */
dout[258]= { 10'sd511   , -10'sd13    }; /* W[   4] =  0.9980  -0.0254i */
dout[259]= { 10'sd511   , -10'sd19    }; /* W[   6] =  0.9980  -0.0371i */
dout[260]= { 10'sd511   , -10'sd25    }; /* W[   8] =  0.9980  -0.0488i */
dout[261]= { 10'sd511   , -10'sd31    }; /* W[  10] =  0.9980  -0.0605i */
dout[262]= { 10'sd511   , -10'sd38    }; /* W[  12] =  0.9980  -0.0742i */
dout[263]= { 10'sd510   , -10'sd44    }; /* W[  14] =  0.9961  -0.0859i */
dout[264]= { 10'sd510   , -10'sd50    }; /* W[  16] =  0.9961  -0.0977i */
dout[265]= { 10'sd509   , -10'sd56    }; /* W[  18] =  0.9941  -0.1094i */
dout[266]= { 10'sd508   , -10'sd63    }; /* W[  20] =  0.9922  -0.1230i */
dout[267]= { 10'sd507   , -10'sd69    }; /* W[  22] =  0.9902  -0.1348i */
dout[268]= { 10'sd506   , -10'sd75    }; /* W[  24] =  0.9883  -0.1465i */
dout[269]= { 10'sd505   , -10'sd81    }; /* W[  26] =  0.9863  -0.1582i */
dout[270]= { 10'sd504   , -10'sd88    }; /* W[  28] =  0.9844  -0.1719i */
dout[271]= { 10'sd503   , -10'sd94    }; /* W[  30] =  0.9824  -0.1836i */
dout[272]= { 10'sd502   , -10'sd100   }; /* W[  32] =  0.9805  -0.1953i */
dout[273]= { 10'sd501   , -10'sd106   }; /* W[  34] =  0.9785  -0.2070i */
dout[274]= { 10'sd500   , -10'sd112   }; /* W[  36] =  0.9766  -0.2188i */
dout[275]= { 10'sd498   , -10'sd118   }; /* W[  38] =  0.9727  -0.2305i */
dout[276]= { 10'sd497   , -10'sd124   }; /* W[  40] =  0.9707  -0.2422i */
dout[277]= { 10'sd495   , -10'sd130   }; /* W[  42] =  0.9668  -0.2539i */
dout[278]= { 10'sd493   , -10'sd137   }; /* W[  44] =  0.9629  -0.2676i */
dout[279]= { 10'sd492   , -10'sd143   }; /* W[  46] =  0.9609  -0.2793i */
dout[280]= { 10'sd490   , -10'sd149   }; /* W[  48] =  0.9570  -0.2910i */
dout[281]= { 10'sd488   , -10'sd155   }; /* W[  50] =  0.9531  -0.3027i */
dout[282]= { 10'sd486   , -10'sd161   }; /* W[  52] =  0.9492  -0.3145i */
dout[283]= { 10'sd484   , -10'sd167   }; /* W[  54] =  0.9453  -0.3262i */
dout[284]= { 10'sd482   , -10'sd172   }; /* W[  56] =  0.9414  -0.3359i */
dout[285]= { 10'sd480   , -10'sd178   }; /* W[  58] =  0.9375  -0.3477i */
dout[286]= { 10'sd478   , -10'sd184   }; /* W[  60] =  0.9336  -0.3594i */
dout[287]= { 10'sd475   , -10'sd190   }; /* W[  62] =  0.9277  -0.3711i */
dout[288]= { 10'sd473   , -10'sd196   }; /* W[  64] =  0.9238  -0.3828i */
dout[289]= { 10'sd471   , -10'sd202   }; /* W[  66] =  0.9199  -0.3945i */
dout[290]= { 10'sd468   , -10'sd207   }; /* W[  68] =  0.9141  -0.4043i */
dout[291]= { 10'sd465   , -10'sd213   }; /* W[  70] =  0.9082  -0.4160i */
dout[292]= { 10'sd463   , -10'sd219   }; /* W[  72] =  0.9043  -0.4277i */
dout[293]= { 10'sd460   , -10'sd225   }; /* W[  74] =  0.8984  -0.4395i */
dout[294]= { 10'sd457   , -10'sd230   }; /* W[  76] =  0.8926  -0.4492i */
dout[295]= { 10'sd454   , -10'sd236   }; /* W[  78] =  0.8867  -0.4609i */
dout[296]= { 10'sd452   , -10'sd241   }; /* W[  80] =  0.8828  -0.4707i */
dout[297]= { 10'sd449   , -10'sd247   }; /* W[  82] =  0.8770  -0.4824i */
dout[298]= { 10'sd445   , -10'sd252   }; /* W[  84] =  0.8691  -0.4922i */
dout[299]= { 10'sd442   , -10'sd258   }; /* W[  86] =  0.8633  -0.5039i */
dout[300]= { 10'sd439   , -10'sd263   }; /* W[  88] =  0.8574  -0.5137i */
dout[301]= { 10'sd436   , -10'sd269   }; /* W[  90] =  0.8516  -0.5254i */
dout[302]= { 10'sd433   , -10'sd274   }; /* W[  92] =  0.8457  -0.5352i */
dout[303]= { 10'sd429   , -10'sd279   }; /* W[  94] =  0.8379  -0.5449i */
dout[304]= { 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[305]= { 10'sd422   , -10'sd290   }; /* W[  98] =  0.8242  -0.5664i */
dout[306]= { 10'sd419   , -10'sd295   }; /* W[ 100] =  0.8184  -0.5762i */
dout[307]= { 10'sd415   , -10'sd300   }; /* W[ 102] =  0.8105  -0.5859i */
dout[308]= { 10'sd411   , -10'sd305   }; /* W[ 104] =  0.8027  -0.5957i */
dout[309]= { 10'sd407   , -10'sd310   }; /* W[ 106] =  0.7949  -0.6055i */
dout[310]= { 10'sd404   , -10'sd315   }; /* W[ 108] =  0.7891  -0.6152i */
dout[311]= { 10'sd400   , -10'sd320   }; /* W[ 110] =  0.7812  -0.6250i */
dout[312]= { 10'sd396   , -10'sd325   }; /* W[ 112] =  0.7734  -0.6348i */
dout[313]= { 10'sd392   , -10'sd330   }; /* W[ 114] =  0.7656  -0.6445i */
dout[314]= { 10'sd388   , -10'sd334   }; /* W[ 116] =  0.7578  -0.6523i */
dout[315]= { 10'sd384   , -10'sd339   }; /* W[ 118] =  0.7500  -0.6621i */
dout[316]= { 10'sd379   , -10'sd344   }; /* W[ 120] =  0.7402  -0.6719i */
dout[317]= { 10'sd375   , -10'sd348   }; /* W[ 122] =  0.7324  -0.6797i */
dout[318]= { 10'sd371   , -10'sd353   }; /* W[ 124] =  0.7246  -0.6895i */
dout[319]= { 10'sd366   , -10'sd358   }; /* W[ 126] =  0.7148  -0.6992i */
dout[320]= { 10'sd362   , -10'sd362   }; /* W[ 128] =  0.7070  -0.7070i */
dout[321]= { 10'sd358   , -10'sd366   }; /* W[ 130] =  0.6992  -0.7148i */
dout[322]= { 10'sd353   , -10'sd371   }; /* W[ 132] =  0.6895  -0.7246i */
dout[323]= { 10'sd348   , -10'sd375   }; /* W[ 134] =  0.6797  -0.7324i */
dout[324]= { 10'sd344   , -10'sd379   }; /* W[ 136] =  0.6719  -0.7402i */
dout[325]= { 10'sd339   , -10'sd384   }; /* W[ 138] =  0.6621  -0.7500i */
dout[326]= { 10'sd334   , -10'sd388   }; /* W[ 140] =  0.6523  -0.7578i */
dout[327]= { 10'sd330   , -10'sd392   }; /* W[ 142] =  0.6445  -0.7656i */
dout[328]= { 10'sd325   , -10'sd396   }; /* W[ 144] =  0.6348  -0.7734i */
dout[329]= { 10'sd320   , -10'sd400   }; /* W[ 146] =  0.6250  -0.7812i */
dout[330]= { 10'sd315   , -10'sd404   }; /* W[ 148] =  0.6152  -0.7891i */
dout[331]= { 10'sd310   , -10'sd407   }; /* W[ 150] =  0.6055  -0.7949i */
dout[332]= { 10'sd305   , -10'sd411   }; /* W[ 152] =  0.5957  -0.8027i */
dout[333]= { 10'sd300   , -10'sd415   }; /* W[ 154] =  0.5859  -0.8105i */
dout[334]= { 10'sd295   , -10'sd419   }; /* W[ 156] =  0.5762  -0.8184i */
dout[335]= { 10'sd290   , -10'sd422   }; /* W[ 158] =  0.5664  -0.8242i */
dout[336]= { 10'sd284   , -10'sd426   }; /* W[ 160] =  0.5547  -0.8320i */
dout[337]= { 10'sd279   , -10'sd429   }; /* W[ 162] =  0.5449  -0.8379i */
dout[338]= { 10'sd274   , -10'sd433   }; /* W[ 164] =  0.5352  -0.8457i */
dout[339]= { 10'sd269   , -10'sd436   }; /* W[ 166] =  0.5254  -0.8516i */
dout[340]= { 10'sd263   , -10'sd439   }; /* W[ 168] =  0.5137  -0.8574i */
dout[341]= { 10'sd258   , -10'sd442   }; /* W[ 170] =  0.5039  -0.8633i */
dout[342]= { 10'sd252   , -10'sd445   }; /* W[ 172] =  0.4922  -0.8691i */
dout[343]= { 10'sd247   , -10'sd449   }; /* W[ 174] =  0.4824  -0.8770i */
dout[344]= { 10'sd241   , -10'sd452   }; /* W[ 176] =  0.4707  -0.8828i */
dout[345]= { 10'sd236   , -10'sd454   }; /* W[ 178] =  0.4609  -0.8867i */
dout[346]= { 10'sd230   , -10'sd457   }; /* W[ 180] =  0.4492  -0.8926i */
dout[347]= { 10'sd225   , -10'sd460   }; /* W[ 182] =  0.4395  -0.8984i */
dout[348]= { 10'sd219   , -10'sd463   }; /* W[ 184] =  0.4277  -0.9043i */
dout[349]= { 10'sd213   , -10'sd465   }; /* W[ 186] =  0.4160  -0.9082i */
dout[350]= { 10'sd207   , -10'sd468   }; /* W[ 188] =  0.4043  -0.9141i */
dout[351]= { 10'sd202   , -10'sd471   }; /* W[ 190] =  0.3945  -0.9199i */
dout[352]= { 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[353]= { 10'sd190   , -10'sd475   }; /* W[ 194] =  0.3711  -0.9277i */
dout[354]= { 10'sd184   , -10'sd478   }; /* W[ 196] =  0.3594  -0.9336i */
dout[355]= { 10'sd178   , -10'sd480   }; /* W[ 198] =  0.3477  -0.9375i */
dout[356]= { 10'sd172   , -10'sd482   }; /* W[ 200] =  0.3359  -0.9414i */
dout[357]= { 10'sd167   , -10'sd484   }; /* W[ 202] =  0.3262  -0.9453i */
dout[358]= { 10'sd161   , -10'sd486   }; /* W[ 204] =  0.3145  -0.9492i */
dout[359]= { 10'sd155   , -10'sd488   }; /* W[ 206] =  0.3027  -0.9531i */
dout[360]= { 10'sd149   , -10'sd490   }; /* W[ 208] =  0.2910  -0.9570i */
dout[361]= { 10'sd143   , -10'sd492   }; /* W[ 210] =  0.2793  -0.9609i */
dout[362]= { 10'sd137   , -10'sd493   }; /* W[ 212] =  0.2676  -0.9629i */
dout[363]= { 10'sd130   , -10'sd495   }; /* W[ 214] =  0.2539  -0.9668i */
dout[364]= { 10'sd124   , -10'sd497   }; /* W[ 216] =  0.2422  -0.9707i */
dout[365]= { 10'sd118   , -10'sd498   }; /* W[ 218] =  0.2305  -0.9727i */
dout[366]= { 10'sd112   , -10'sd500   }; /* W[ 220] =  0.2188  -0.9766i */
dout[367]= { 10'sd106   , -10'sd501   }; /* W[ 222] =  0.2070  -0.9785i */
dout[368]= { 10'sd100   , -10'sd502   }; /* W[ 224] =  0.1953  -0.9805i */
dout[369]= { 10'sd94    , -10'sd503   }; /* W[ 226] =  0.1836  -0.9824i */
dout[370]= { 10'sd88    , -10'sd504   }; /* W[ 228] =  0.1719  -0.9844i */
dout[371]= { 10'sd81    , -10'sd505   }; /* W[ 230] =  0.1582  -0.9863i */
dout[372]= { 10'sd75    , -10'sd506   }; /* W[ 232] =  0.1465  -0.9883i */
dout[373]= { 10'sd69    , -10'sd507   }; /* W[ 234] =  0.1348  -0.9902i */
dout[374]= { 10'sd63    , -10'sd508   }; /* W[ 236] =  0.1230  -0.9922i */
dout[375]= { 10'sd56    , -10'sd509   }; /* W[ 238] =  0.1094  -0.9941i */
dout[376]= { 10'sd50    , -10'sd510   }; /* W[ 240] =  0.0977  -0.9961i */
dout[377]= { 10'sd44    , -10'sd510   }; /* W[ 242] =  0.0859  -0.9961i */
dout[378]= { 10'sd38    , -10'sd511   }; /* W[ 244] =  0.0742  -0.9980i */
dout[379]= { 10'sd31    , -10'sd511   }; /* W[ 246] =  0.0605  -0.9980i */
dout[380]= { 10'sd25    , -10'sd511   }; /* W[ 248] =  0.0488  -0.9980i */
dout[381]= { 10'sd19    , -10'sd512   }; /* W[ 250] =  0.0371  -1.0000i */
dout[382]= { 10'sd13    , -10'sd512   }; /* W[ 252] =  0.0254  -1.0000i */
dout[383]= { 10'sd6     , -10'sd512   }; /* W[ 254] =  0.0117  -1.0000i */
dout[384]= { 10'sd0     , -10'sd512   }; /* W[ 256] =  0.0000  -1.0000i */
dout[385]= {-10'sd6     , -10'sd512   }; /* W[ 258] = -0.0117  -1.0000i */
dout[386]= {-10'sd13    , -10'sd512   }; /* W[ 260] = -0.0254  -1.0000i */
dout[387]= {-10'sd19    , -10'sd512   }; /* W[ 262] = -0.0371  -1.0000i */
dout[388]= {-10'sd25    , -10'sd511   }; /* W[ 264] = -0.0488  -0.9980i */
dout[389]= {-10'sd31    , -10'sd511   }; /* W[ 266] = -0.0605  -0.9980i */
dout[390]= {-10'sd38    , -10'sd511   }; /* W[ 268] = -0.0742  -0.9980i */
dout[391]= {-10'sd44    , -10'sd510   }; /* W[ 270] = -0.0859  -0.9961i */
dout[392]= {-10'sd50    , -10'sd510   }; /* W[ 272] = -0.0977  -0.9961i */
dout[393]= {-10'sd56    , -10'sd509   }; /* W[ 274] = -0.1094  -0.9941i */
dout[394]= {-10'sd63    , -10'sd508   }; /* W[ 276] = -0.1230  -0.9922i */
dout[395]= {-10'sd69    , -10'sd507   }; /* W[ 278] = -0.1348  -0.9902i */
dout[396]= {-10'sd75    , -10'sd506   }; /* W[ 280] = -0.1465  -0.9883i */
dout[397]= {-10'sd81    , -10'sd505   }; /* W[ 282] = -0.1582  -0.9863i */
dout[398]= {-10'sd88    , -10'sd504   }; /* W[ 284] = -0.1719  -0.9844i */
dout[399]= {-10'sd94    , -10'sd503   }; /* W[ 286] = -0.1836  -0.9824i */
dout[400]= {-10'sd100   , -10'sd502   }; /* W[ 288] = -0.1953  -0.9805i */
dout[401]= {-10'sd106   , -10'sd501   }; /* W[ 290] = -0.2070  -0.9785i */
dout[402]= {-10'sd112   , -10'sd500   }; /* W[ 292] = -0.2188  -0.9766i */
dout[403]= {-10'sd118   , -10'sd498   }; /* W[ 294] = -0.2305  -0.9727i */
dout[404]= {-10'sd124   , -10'sd497   }; /* W[ 296] = -0.2422  -0.9707i */
dout[405]= {-10'sd130   , -10'sd495   }; /* W[ 298] = -0.2539  -0.9668i */
dout[406]= {-10'sd137   , -10'sd493   }; /* W[ 300] = -0.2676  -0.9629i */
dout[407]= {-10'sd143   , -10'sd492   }; /* W[ 302] = -0.2793  -0.9609i */
dout[408]= {-10'sd149   , -10'sd490   }; /* W[ 304] = -0.2910  -0.9570i */
dout[409]= {-10'sd155   , -10'sd488   }; /* W[ 306] = -0.3027  -0.9531i */
dout[410]= {-10'sd161   , -10'sd486   }; /* W[ 308] = -0.3145  -0.9492i */
dout[411]= {-10'sd167   , -10'sd484   }; /* W[ 310] = -0.3262  -0.9453i */
dout[412]= {-10'sd172   , -10'sd482   }; /* W[ 312] = -0.3359  -0.9414i */
dout[413]= {-10'sd178   , -10'sd480   }; /* W[ 314] = -0.3477  -0.9375i */
dout[414]= {-10'sd184   , -10'sd478   }; /* W[ 316] = -0.3594  -0.9336i */
dout[415]= {-10'sd190   , -10'sd475   }; /* W[ 318] = -0.3711  -0.9277i */
dout[416]= {-10'sd196   , -10'sd473   }; /* W[ 320] = -0.3828  -0.9238i */
dout[417]= {-10'sd202   , -10'sd471   }; /* W[ 322] = -0.3945  -0.9199i */
dout[418]= {-10'sd207   , -10'sd468   }; /* W[ 324] = -0.4043  -0.9141i */
dout[419]= {-10'sd213   , -10'sd465   }; /* W[ 326] = -0.4160  -0.9082i */
dout[420]= {-10'sd219   , -10'sd463   }; /* W[ 328] = -0.4277  -0.9043i */
dout[421]= {-10'sd225   , -10'sd460   }; /* W[ 330] = -0.4395  -0.8984i */
dout[422]= {-10'sd230   , -10'sd457   }; /* W[ 332] = -0.4492  -0.8926i */
dout[423]= {-10'sd236   , -10'sd454   }; /* W[ 334] = -0.4609  -0.8867i */
dout[424]= {-10'sd241   , -10'sd452   }; /* W[ 336] = -0.4707  -0.8828i */
dout[425]= {-10'sd247   , -10'sd449   }; /* W[ 338] = -0.4824  -0.8770i */
dout[426]= {-10'sd252   , -10'sd445   }; /* W[ 340] = -0.4922  -0.8691i */
dout[427]= {-10'sd258   , -10'sd442   }; /* W[ 342] = -0.5039  -0.8633i */
dout[428]= {-10'sd263   , -10'sd439   }; /* W[ 344] = -0.5137  -0.8574i */
dout[429]= {-10'sd269   , -10'sd436   }; /* W[ 346] = -0.5254  -0.8516i */
dout[430]= {-10'sd274   , -10'sd433   }; /* W[ 348] = -0.5352  -0.8457i */
dout[431]= {-10'sd279   , -10'sd429   }; /* W[ 350] = -0.5449  -0.8379i */
dout[432]= {-10'sd284   , -10'sd426   }; /* W[ 352] = -0.5547  -0.8320i */
dout[433]= {-10'sd290   , -10'sd422   }; /* W[ 354] = -0.5664  -0.8242i */
dout[434]= {-10'sd295   , -10'sd419   }; /* W[ 356] = -0.5762  -0.8184i */
dout[435]= {-10'sd300   , -10'sd415   }; /* W[ 358] = -0.5859  -0.8105i */
dout[436]= {-10'sd305   , -10'sd411   }; /* W[ 360] = -0.5957  -0.8027i */
dout[437]= {-10'sd310   , -10'sd407   }; /* W[ 362] = -0.6055  -0.7949i */
dout[438]= {-10'sd315   , -10'sd404   }; /* W[ 364] = -0.6152  -0.7891i */
dout[439]= {-10'sd320   , -10'sd400   }; /* W[ 366] = -0.6250  -0.7812i */
dout[440]= {-10'sd325   , -10'sd396   }; /* W[ 368] = -0.6348  -0.7734i */
dout[441]= {-10'sd330   , -10'sd392   }; /* W[ 370] = -0.6445  -0.7656i */
dout[442]= {-10'sd334   , -10'sd388   }; /* W[ 372] = -0.6523  -0.7578i */
dout[443]= {-10'sd339   , -10'sd384   }; /* W[ 374] = -0.6621  -0.7500i */
dout[444]= {-10'sd344   , -10'sd379   }; /* W[ 376] = -0.6719  -0.7402i */
dout[445]= {-10'sd348   , -10'sd375   }; /* W[ 378] = -0.6797  -0.7324i */
dout[446]= {-10'sd353   , -10'sd371   }; /* W[ 380] = -0.6895  -0.7246i */
dout[447]= {-10'sd358   , -10'sd366   }; /* W[ 382] = -0.6992  -0.7148i */
dout[448]= {-10'sd362   , -10'sd362   }; /* W[ 384] = -0.7070  -0.7070i */
dout[449]= {-10'sd366   , -10'sd358   }; /* W[ 386] = -0.7148  -0.6992i */
dout[450]= {-10'sd371   , -10'sd353   }; /* W[ 388] = -0.7246  -0.6895i */
dout[451]= {-10'sd375   , -10'sd348   }; /* W[ 390] = -0.7324  -0.6797i */
dout[452]= {-10'sd379   , -10'sd344   }; /* W[ 392] = -0.7402  -0.6719i */
dout[453]= {-10'sd384   , -10'sd339   }; /* W[ 394] = -0.7500  -0.6621i */
dout[454]= {-10'sd388   , -10'sd334   }; /* W[ 396] = -0.7578  -0.6523i */
dout[455]= {-10'sd392   , -10'sd330   }; /* W[ 398] = -0.7656  -0.6445i */
dout[456]= {-10'sd396   , -10'sd325   }; /* W[ 400] = -0.7734  -0.6348i */
dout[457]= {-10'sd400   , -10'sd320   }; /* W[ 402] = -0.7812  -0.6250i */
dout[458]= {-10'sd404   , -10'sd315   }; /* W[ 404] = -0.7891  -0.6152i */
dout[459]= {-10'sd407   , -10'sd310   }; /* W[ 406] = -0.7949  -0.6055i */
dout[460]= {-10'sd411   , -10'sd305   }; /* W[ 408] = -0.8027  -0.5957i */
dout[461]= {-10'sd415   , -10'sd300   }; /* W[ 410] = -0.8105  -0.5859i */
dout[462]= {-10'sd419   , -10'sd295   }; /* W[ 412] = -0.8184  -0.5762i */
dout[463]= {-10'sd422   , -10'sd290   }; /* W[ 414] = -0.8242  -0.5664i */
dout[464]= {-10'sd426   , -10'sd284   }; /* W[ 416] = -0.8320  -0.5547i */
dout[465]= {-10'sd429   , -10'sd279   }; /* W[ 418] = -0.8379  -0.5449i */
dout[466]= {-10'sd433   , -10'sd274   }; /* W[ 420] = -0.8457  -0.5352i */
dout[467]= {-10'sd436   , -10'sd269   }; /* W[ 422] = -0.8516  -0.5254i */
dout[468]= {-10'sd439   , -10'sd263   }; /* W[ 424] = -0.8574  -0.5137i */
dout[469]= {-10'sd442   , -10'sd258   }; /* W[ 426] = -0.8633  -0.5039i */
dout[470]= {-10'sd445   , -10'sd252   }; /* W[ 428] = -0.8691  -0.4922i */
dout[471]= {-10'sd449   , -10'sd247   }; /* W[ 430] = -0.8770  -0.4824i */
dout[472]= {-10'sd452   , -10'sd241   }; /* W[ 432] = -0.8828  -0.4707i */
dout[473]= {-10'sd454   , -10'sd236   }; /* W[ 434] = -0.8867  -0.4609i */
dout[474]= {-10'sd457   , -10'sd230   }; /* W[ 436] = -0.8926  -0.4492i */
dout[475]= {-10'sd460   , -10'sd225   }; /* W[ 438] = -0.8984  -0.4395i */
dout[476]= {-10'sd463   , -10'sd219   }; /* W[ 440] = -0.9043  -0.4277i */
dout[477]= {-10'sd465   , -10'sd213   }; /* W[ 442] = -0.9082  -0.4160i */
dout[478]= {-10'sd468   , -10'sd207   }; /* W[ 444] = -0.9141  -0.4043i */
dout[479]= {-10'sd471   , -10'sd202   }; /* W[ 446] = -0.9199  -0.3945i */
dout[480]= {-10'sd473   , -10'sd196   }; /* W[ 448] = -0.9238  -0.3828i */
dout[481]= {-10'sd475   , -10'sd190   }; /* W[ 450] = -0.9277  -0.3711i */
dout[482]= {-10'sd478   , -10'sd184   }; /* W[ 452] = -0.9336  -0.3594i */
dout[483]= {-10'sd480   , -10'sd178   }; /* W[ 454] = -0.9375  -0.3477i */
dout[484]= {-10'sd482   , -10'sd172   }; /* W[ 456] = -0.9414  -0.3359i */
dout[485]= {-10'sd484   , -10'sd167   }; /* W[ 458] = -0.9453  -0.3262i */
dout[486]= {-10'sd486   , -10'sd161   }; /* W[ 460] = -0.9492  -0.3145i */
dout[487]= {-10'sd488   , -10'sd155   }; /* W[ 462] = -0.9531  -0.3027i */
dout[488]= {-10'sd490   , -10'sd149   }; /* W[ 464] = -0.9570  -0.2910i */
dout[489]= {-10'sd492   , -10'sd143   }; /* W[ 466] = -0.9609  -0.2793i */
dout[490]= {-10'sd493   , -10'sd137   }; /* W[ 468] = -0.9629  -0.2676i */
dout[491]= {-10'sd495   , -10'sd130   }; /* W[ 470] = -0.9668  -0.2539i */
dout[492]= {-10'sd497   , -10'sd124   }; /* W[ 472] = -0.9707  -0.2422i */
dout[493]= {-10'sd498   , -10'sd118   }; /* W[ 474] = -0.9727  -0.2305i */
dout[494]= {-10'sd500   , -10'sd112   }; /* W[ 476] = -0.9766  -0.2188i */
dout[495]= {-10'sd501   , -10'sd106   }; /* W[ 478] = -0.9785  -0.2070i */
dout[496]= {-10'sd502   , -10'sd100   }; /* W[ 480] = -0.9805  -0.1953i */
dout[497]= {-10'sd503   , -10'sd94    }; /* W[ 482] = -0.9824  -0.1836i */
dout[498]= {-10'sd504   , -10'sd88    }; /* W[ 484] = -0.9844  -0.1719i */
dout[499]= {-10'sd505   , -10'sd81    }; /* W[ 486] = -0.9863  -0.1582i */
dout[500]= {-10'sd506   , -10'sd75    }; /* W[ 488] = -0.9883  -0.1465i */
dout[501]= {-10'sd507   , -10'sd69    }; /* W[ 490] = -0.9902  -0.1348i */
dout[502]= {-10'sd508   , -10'sd63    }; /* W[ 492] = -0.9922  -0.1230i */
dout[503]= {-10'sd509   , -10'sd56    }; /* W[ 494] = -0.9941  -0.1094i */
dout[504]= {-10'sd510   , -10'sd50    }; /* W[ 496] = -0.9961  -0.0977i */
dout[505]= {-10'sd510   , -10'sd44    }; /* W[ 498] = -0.9961  -0.0859i */
dout[506]= {-10'sd511   , -10'sd38    }; /* W[ 500] = -0.9980  -0.0742i */
dout[507]= {-10'sd511   , -10'sd31    }; /* W[ 502] = -0.9980  -0.0605i */
dout[508]= {-10'sd511   , -10'sd25    }; /* W[ 504] = -0.9980  -0.0488i */
dout[509]= {-10'sd512   , -10'sd19    }; /* W[ 506] = -1.0000  -0.0371i */
dout[510]= {-10'sd512   , -10'sd13    }; /* W[ 508] = -1.0000  -0.0254i */
dout[511]= {-10'sd512   , -10'sd6     }; /* W[ 510] = -1.0000  -0.0117i */
dout[512]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[513]= { 10'sd511   , -10'sd3     }; /* W[   1] =  0.9980  -0.0059i */
dout[514]= { 10'sd511   , -10'sd6     }; /* W[   2] =  0.9980  -0.0117i */
dout[515]= { 10'sd511   , -10'sd9     }; /* W[   3] =  0.9980  -0.0176i */
dout[516]= { 10'sd511   , -10'sd13    }; /* W[   4] =  0.9980  -0.0254i */
dout[517]= { 10'sd511   , -10'sd16    }; /* W[   5] =  0.9980  -0.0312i */
dout[518]= { 10'sd511   , -10'sd19    }; /* W[   6] =  0.9980  -0.0371i */
dout[519]= { 10'sd511   , -10'sd22    }; /* W[   7] =  0.9980  -0.0430i */
dout[520]= { 10'sd511   , -10'sd25    }; /* W[   8] =  0.9980  -0.0488i */
dout[521]= { 10'sd511   , -10'sd28    }; /* W[   9] =  0.9980  -0.0547i */
dout[522]= { 10'sd511   , -10'sd31    }; /* W[  10] =  0.9980  -0.0605i */
dout[523]= { 10'sd511   , -10'sd35    }; /* W[  11] =  0.9980  -0.0684i */
dout[524]= { 10'sd511   , -10'sd38    }; /* W[  12] =  0.9980  -0.0742i */
dout[525]= { 10'sd510   , -10'sd41    }; /* W[  13] =  0.9961  -0.0801i */
dout[526]= { 10'sd510   , -10'sd44    }; /* W[  14] =  0.9961  -0.0859i */
dout[527]= { 10'sd510   , -10'sd47    }; /* W[  15] =  0.9961  -0.0918i */
dout[528]= { 10'sd510   , -10'sd50    }; /* W[  16] =  0.9961  -0.0977i */
dout[529]= { 10'sd509   , -10'sd53    }; /* W[  17] =  0.9941  -0.1035i */
dout[530]= { 10'sd509   , -10'sd56    }; /* W[  18] =  0.9941  -0.1094i */
dout[531]= { 10'sd509   , -10'sd60    }; /* W[  19] =  0.9941  -0.1172i */
dout[532]= { 10'sd508   , -10'sd63    }; /* W[  20] =  0.9922  -0.1230i */
dout[533]= { 10'sd508   , -10'sd66    }; /* W[  21] =  0.9922  -0.1289i */
dout[534]= { 10'sd507   , -10'sd69    }; /* W[  22] =  0.9902  -0.1348i */
dout[535]= { 10'sd507   , -10'sd72    }; /* W[  23] =  0.9902  -0.1406i */
dout[536]= { 10'sd506   , -10'sd75    }; /* W[  24] =  0.9883  -0.1465i */
dout[537]= { 10'sd506   , -10'sd78    }; /* W[  25] =  0.9883  -0.1523i */
dout[538]= { 10'sd505   , -10'sd81    }; /* W[  26] =  0.9863  -0.1582i */
dout[539]= { 10'sd505   , -10'sd84    }; /* W[  27] =  0.9863  -0.1641i */
dout[540]= { 10'sd504   , -10'sd88    }; /* W[  28] =  0.9844  -0.1719i */
dout[541]= { 10'sd504   , -10'sd91    }; /* W[  29] =  0.9844  -0.1777i */
dout[542]= { 10'sd503   , -10'sd94    }; /* W[  30] =  0.9824  -0.1836i */
dout[543]= { 10'sd503   , -10'sd97    }; /* W[  31] =  0.9824  -0.1895i */
dout[544]= { 10'sd502   , -10'sd100   }; /* W[  32] =  0.9805  -0.1953i */
dout[545]= { 10'sd502   , -10'sd103   }; /* W[  33] =  0.9805  -0.2012i */
dout[546]= { 10'sd501   , -10'sd106   }; /* W[  34] =  0.9785  -0.2070i */
dout[547]= { 10'sd500   , -10'sd109   }; /* W[  35] =  0.9766  -0.2129i */
dout[548]= { 10'sd500   , -10'sd112   }; /* W[  36] =  0.9766  -0.2188i */
dout[549]= { 10'sd499   , -10'sd115   }; /* W[  37] =  0.9746  -0.2246i */
dout[550]= { 10'sd498   , -10'sd118   }; /* W[  38] =  0.9727  -0.2305i */
dout[551]= { 10'sd497   , -10'sd121   }; /* W[  39] =  0.9707  -0.2363i */
dout[552]= { 10'sd497   , -10'sd124   }; /* W[  40] =  0.9707  -0.2422i */
dout[553]= { 10'sd496   , -10'sd127   }; /* W[  41] =  0.9688  -0.2480i */
dout[554]= { 10'sd495   , -10'sd130   }; /* W[  42] =  0.9668  -0.2539i */
dout[555]= { 10'sd494   , -10'sd134   }; /* W[  43] =  0.9648  -0.2617i */
dout[556]= { 10'sd493   , -10'sd137   }; /* W[  44] =  0.9629  -0.2676i */
dout[557]= { 10'sd493   , -10'sd140   }; /* W[  45] =  0.9629  -0.2734i */
dout[558]= { 10'sd492   , -10'sd143   }; /* W[  46] =  0.9609  -0.2793i */
dout[559]= { 10'sd491   , -10'sd146   }; /* W[  47] =  0.9590  -0.2852i */
dout[560]= { 10'sd490   , -10'sd149   }; /* W[  48] =  0.9570  -0.2910i */
dout[561]= { 10'sd489   , -10'sd152   }; /* W[  49] =  0.9551  -0.2969i */
dout[562]= { 10'sd488   , -10'sd155   }; /* W[  50] =  0.9531  -0.3027i */
dout[563]= { 10'sd487   , -10'sd158   }; /* W[  51] =  0.9512  -0.3086i */
dout[564]= { 10'sd486   , -10'sd161   }; /* W[  52] =  0.9492  -0.3145i */
dout[565]= { 10'sd485   , -10'sd164   }; /* W[  53] =  0.9473  -0.3203i */
dout[566]= { 10'sd484   , -10'sd167   }; /* W[  54] =  0.9453  -0.3262i */
dout[567]= { 10'sd483   , -10'sd170   }; /* W[  55] =  0.9434  -0.3320i */
dout[568]= { 10'sd482   , -10'sd172   }; /* W[  56] =  0.9414  -0.3359i */
dout[569]= { 10'sd481   , -10'sd175   }; /* W[  57] =  0.9395  -0.3418i */
dout[570]= { 10'sd480   , -10'sd178   }; /* W[  58] =  0.9375  -0.3477i */
dout[571]= { 10'sd479   , -10'sd181   }; /* W[  59] =  0.9355  -0.3535i */
dout[572]= { 10'sd478   , -10'sd184   }; /* W[  60] =  0.9336  -0.3594i */
dout[573]= { 10'sd477   , -10'sd187   }; /* W[  61] =  0.9316  -0.3652i */
dout[574]= { 10'sd475   , -10'sd190   }; /* W[  62] =  0.9277  -0.3711i */
dout[575]= { 10'sd474   , -10'sd193   }; /* W[  63] =  0.9258  -0.3770i */
dout[576]= { 10'sd473   , -10'sd196   }; /* W[  64] =  0.9238  -0.3828i */
dout[577]= { 10'sd472   , -10'sd199   }; /* W[  65] =  0.9219  -0.3887i */
dout[578]= { 10'sd471   , -10'sd202   }; /* W[  66] =  0.9199  -0.3945i */
dout[579]= { 10'sd469   , -10'sd205   }; /* W[  67] =  0.9160  -0.4004i */
dout[580]= { 10'sd468   , -10'sd207   }; /* W[  68] =  0.9141  -0.4043i */
dout[581]= { 10'sd467   , -10'sd210   }; /* W[  69] =  0.9121  -0.4102i */
dout[582]= { 10'sd465   , -10'sd213   }; /* W[  70] =  0.9082  -0.4160i */
dout[583]= { 10'sd464   , -10'sd216   }; /* W[  71] =  0.9062  -0.4219i */
dout[584]= { 10'sd463   , -10'sd219   }; /* W[  72] =  0.9043  -0.4277i */
dout[585]= { 10'sd461   , -10'sd222   }; /* W[  73] =  0.9004  -0.4336i */
dout[586]= { 10'sd460   , -10'sd225   }; /* W[  74] =  0.8984  -0.4395i */
dout[587]= { 10'sd459   , -10'sd227   }; /* W[  75] =  0.8965  -0.4434i */
dout[588]= { 10'sd457   , -10'sd230   }; /* W[  76] =  0.8926  -0.4492i */
dout[589]= { 10'sd456   , -10'sd233   }; /* W[  77] =  0.8906  -0.4551i */
dout[590]= { 10'sd454   , -10'sd236   }; /* W[  78] =  0.8867  -0.4609i */
dout[591]= { 10'sd453   , -10'sd239   }; /* W[  79] =  0.8848  -0.4668i */
dout[592]= { 10'sd452   , -10'sd241   }; /* W[  80] =  0.8828  -0.4707i */
dout[593]= { 10'sd450   , -10'sd244   }; /* W[  81] =  0.8789  -0.4766i */
dout[594]= { 10'sd449   , -10'sd247   }; /* W[  82] =  0.8770  -0.4824i */
dout[595]= { 10'sd447   , -10'sd250   }; /* W[  83] =  0.8730  -0.4883i */
dout[596]= { 10'sd445   , -10'sd252   }; /* W[  84] =  0.8691  -0.4922i */
dout[597]= { 10'sd444   , -10'sd255   }; /* W[  85] =  0.8672  -0.4980i */
dout[598]= { 10'sd442   , -10'sd258   }; /* W[  86] =  0.8633  -0.5039i */
dout[599]= { 10'sd441   , -10'sd261   }; /* W[  87] =  0.8613  -0.5098i */
dout[600]= { 10'sd439   , -10'sd263   }; /* W[  88] =  0.8574  -0.5137i */
dout[601]= { 10'sd438   , -10'sd266   }; /* W[  89] =  0.8555  -0.5195i */
dout[602]= { 10'sd436   , -10'sd269   }; /* W[  90] =  0.8516  -0.5254i */
dout[603]= { 10'sd434   , -10'sd271   }; /* W[  91] =  0.8477  -0.5293i */
dout[604]= { 10'sd433   , -10'sd274   }; /* W[  92] =  0.8457  -0.5352i */
dout[605]= { 10'sd431   , -10'sd277   }; /* W[  93] =  0.8418  -0.5410i */
dout[606]= { 10'sd429   , -10'sd279   }; /* W[  94] =  0.8379  -0.5449i */
dout[607]= { 10'sd427   , -10'sd282   }; /* W[  95] =  0.8340  -0.5508i */
dout[608]= { 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[609]= { 10'sd424   , -10'sd287   }; /* W[  97] =  0.8281  -0.5605i */
dout[610]= { 10'sd422   , -10'sd290   }; /* W[  98] =  0.8242  -0.5664i */
dout[611]= { 10'sd420   , -10'sd292   }; /* W[  99] =  0.8203  -0.5703i */
dout[612]= { 10'sd419   , -10'sd295   }; /* W[ 100] =  0.8184  -0.5762i */
dout[613]= { 10'sd417   , -10'sd297   }; /* W[ 101] =  0.8145  -0.5801i */
dout[614]= { 10'sd415   , -10'sd300   }; /* W[ 102] =  0.8105  -0.5859i */
dout[615]= { 10'sd413   , -10'sd302   }; /* W[ 103] =  0.8066  -0.5898i */
dout[616]= { 10'sd411   , -10'sd305   }; /* W[ 104] =  0.8027  -0.5957i */
dout[617]= { 10'sd409   , -10'sd308   }; /* W[ 105] =  0.7988  -0.6016i */
dout[618]= { 10'sd407   , -10'sd310   }; /* W[ 106] =  0.7949  -0.6055i */
dout[619]= { 10'sd406   , -10'sd313   }; /* W[ 107] =  0.7930  -0.6113i */
dout[620]= { 10'sd404   , -10'sd315   }; /* W[ 108] =  0.7891  -0.6152i */
dout[621]= { 10'sd402   , -10'sd317   }; /* W[ 109] =  0.7852  -0.6191i */
dout[622]= { 10'sd400   , -10'sd320   }; /* W[ 110] =  0.7812  -0.6250i */
dout[623]= { 10'sd398   , -10'sd322   }; /* W[ 111] =  0.7773  -0.6289i */
dout[624]= { 10'sd396   , -10'sd325   }; /* W[ 112] =  0.7734  -0.6348i */
dout[625]= { 10'sd394   , -10'sd327   }; /* W[ 113] =  0.7695  -0.6387i */
dout[626]= { 10'sd392   , -10'sd330   }; /* W[ 114] =  0.7656  -0.6445i */
dout[627]= { 10'sd390   , -10'sd332   }; /* W[ 115] =  0.7617  -0.6484i */
dout[628]= { 10'sd388   , -10'sd334   }; /* W[ 116] =  0.7578  -0.6523i */
dout[629]= { 10'sd386   , -10'sd337   }; /* W[ 117] =  0.7539  -0.6582i */
dout[630]= { 10'sd384   , -10'sd339   }; /* W[ 118] =  0.7500  -0.6621i */
dout[631]= { 10'sd381   , -10'sd342   }; /* W[ 119] =  0.7441  -0.6680i */
dout[632]= { 10'sd379   , -10'sd344   }; /* W[ 120] =  0.7402  -0.6719i */
dout[633]= { 10'sd377   , -10'sd346   }; /* W[ 121] =  0.7363  -0.6758i */
dout[634]= { 10'sd375   , -10'sd348   }; /* W[ 122] =  0.7324  -0.6797i */
dout[635]= { 10'sd373   , -10'sd351   }; /* W[ 123] =  0.7285  -0.6855i */
dout[636]= { 10'sd371   , -10'sd353   }; /* W[ 124] =  0.7246  -0.6895i */
dout[637]= { 10'sd369   , -10'sd355   }; /* W[ 125] =  0.7207  -0.6934i */
dout[638]= { 10'sd366   , -10'sd358   }; /* W[ 126] =  0.7148  -0.6992i */
dout[639]= { 10'sd364   , -10'sd360   }; /* W[ 127] =  0.7109  -0.7031i */
dout[640]= { 10'sd362   , -10'sd362   }; /* W[ 128] =  0.7070  -0.7070i */
dout[641]= { 10'sd360   , -10'sd364   }; /* W[ 129] =  0.7031  -0.7109i */
dout[642]= { 10'sd358   , -10'sd366   }; /* W[ 130] =  0.6992  -0.7148i */
dout[643]= { 10'sd355   , -10'sd369   }; /* W[ 131] =  0.6934  -0.7207i */
dout[644]= { 10'sd353   , -10'sd371   }; /* W[ 132] =  0.6895  -0.7246i */
dout[645]= { 10'sd351   , -10'sd373   }; /* W[ 133] =  0.6855  -0.7285i */
dout[646]= { 10'sd348   , -10'sd375   }; /* W[ 134] =  0.6797  -0.7324i */
dout[647]= { 10'sd346   , -10'sd377   }; /* W[ 135] =  0.6758  -0.7363i */
dout[648]= { 10'sd344   , -10'sd379   }; /* W[ 136] =  0.6719  -0.7402i */
dout[649]= { 10'sd342   , -10'sd381   }; /* W[ 137] =  0.6680  -0.7441i */
dout[650]= { 10'sd339   , -10'sd384   }; /* W[ 138] =  0.6621  -0.7500i */
dout[651]= { 10'sd337   , -10'sd386   }; /* W[ 139] =  0.6582  -0.7539i */
dout[652]= { 10'sd334   , -10'sd388   }; /* W[ 140] =  0.6523  -0.7578i */
dout[653]= { 10'sd332   , -10'sd390   }; /* W[ 141] =  0.6484  -0.7617i */
dout[654]= { 10'sd330   , -10'sd392   }; /* W[ 142] =  0.6445  -0.7656i */
dout[655]= { 10'sd327   , -10'sd394   }; /* W[ 143] =  0.6387  -0.7695i */
dout[656]= { 10'sd325   , -10'sd396   }; /* W[ 144] =  0.6348  -0.7734i */
dout[657]= { 10'sd322   , -10'sd398   }; /* W[ 145] =  0.6289  -0.7773i */
dout[658]= { 10'sd320   , -10'sd400   }; /* W[ 146] =  0.6250  -0.7812i */
dout[659]= { 10'sd317   , -10'sd402   }; /* W[ 147] =  0.6191  -0.7852i */
dout[660]= { 10'sd315   , -10'sd404   }; /* W[ 148] =  0.6152  -0.7891i */
dout[661]= { 10'sd313   , -10'sd406   }; /* W[ 149] =  0.6113  -0.7930i */
dout[662]= { 10'sd310   , -10'sd407   }; /* W[ 150] =  0.6055  -0.7949i */
dout[663]= { 10'sd308   , -10'sd409   }; /* W[ 151] =  0.6016  -0.7988i */
dout[664]= { 10'sd305   , -10'sd411   }; /* W[ 152] =  0.5957  -0.8027i */
dout[665]= { 10'sd302   , -10'sd413   }; /* W[ 153] =  0.5898  -0.8066i */
dout[666]= { 10'sd300   , -10'sd415   }; /* W[ 154] =  0.5859  -0.8105i */
dout[667]= { 10'sd297   , -10'sd417   }; /* W[ 155] =  0.5801  -0.8145i */
dout[668]= { 10'sd295   , -10'sd419   }; /* W[ 156] =  0.5762  -0.8184i */
dout[669]= { 10'sd292   , -10'sd420   }; /* W[ 157] =  0.5703  -0.8203i */
dout[670]= { 10'sd290   , -10'sd422   }; /* W[ 158] =  0.5664  -0.8242i */
dout[671]= { 10'sd287   , -10'sd424   }; /* W[ 159] =  0.5605  -0.8281i */
dout[672]= { 10'sd284   , -10'sd426   }; /* W[ 160] =  0.5547  -0.8320i */
dout[673]= { 10'sd282   , -10'sd427   }; /* W[ 161] =  0.5508  -0.8340i */
dout[674]= { 10'sd279   , -10'sd429   }; /* W[ 162] =  0.5449  -0.8379i */
dout[675]= { 10'sd277   , -10'sd431   }; /* W[ 163] =  0.5410  -0.8418i */
dout[676]= { 10'sd274   , -10'sd433   }; /* W[ 164] =  0.5352  -0.8457i */
dout[677]= { 10'sd271   , -10'sd434   }; /* W[ 165] =  0.5293  -0.8477i */
dout[678]= { 10'sd269   , -10'sd436   }; /* W[ 166] =  0.5254  -0.8516i */
dout[679]= { 10'sd266   , -10'sd438   }; /* W[ 167] =  0.5195  -0.8555i */
dout[680]= { 10'sd263   , -10'sd439   }; /* W[ 168] =  0.5137  -0.8574i */
dout[681]= { 10'sd261   , -10'sd441   }; /* W[ 169] =  0.5098  -0.8613i */
dout[682]= { 10'sd258   , -10'sd442   }; /* W[ 170] =  0.5039  -0.8633i */
dout[683]= { 10'sd255   , -10'sd444   }; /* W[ 171] =  0.4980  -0.8672i */
dout[684]= { 10'sd252   , -10'sd445   }; /* W[ 172] =  0.4922  -0.8691i */
dout[685]= { 10'sd250   , -10'sd447   }; /* W[ 173] =  0.4883  -0.8730i */
dout[686]= { 10'sd247   , -10'sd449   }; /* W[ 174] =  0.4824  -0.8770i */
dout[687]= { 10'sd244   , -10'sd450   }; /* W[ 175] =  0.4766  -0.8789i */
dout[688]= { 10'sd241   , -10'sd452   }; /* W[ 176] =  0.4707  -0.8828i */
dout[689]= { 10'sd239   , -10'sd453   }; /* W[ 177] =  0.4668  -0.8848i */
dout[690]= { 10'sd236   , -10'sd454   }; /* W[ 178] =  0.4609  -0.8867i */
dout[691]= { 10'sd233   , -10'sd456   }; /* W[ 179] =  0.4551  -0.8906i */
dout[692]= { 10'sd230   , -10'sd457   }; /* W[ 180] =  0.4492  -0.8926i */
dout[693]= { 10'sd227   , -10'sd459   }; /* W[ 181] =  0.4434  -0.8965i */
dout[694]= { 10'sd225   , -10'sd460   }; /* W[ 182] =  0.4395  -0.8984i */
dout[695]= { 10'sd222   , -10'sd461   }; /* W[ 183] =  0.4336  -0.9004i */
dout[696]= { 10'sd219   , -10'sd463   }; /* W[ 184] =  0.4277  -0.9043i */
dout[697]= { 10'sd216   , -10'sd464   }; /* W[ 185] =  0.4219  -0.9062i */
dout[698]= { 10'sd213   , -10'sd465   }; /* W[ 186] =  0.4160  -0.9082i */
dout[699]= { 10'sd210   , -10'sd467   }; /* W[ 187] =  0.4102  -0.9121i */
dout[700]= { 10'sd207   , -10'sd468   }; /* W[ 188] =  0.4043  -0.9141i */
dout[701]= { 10'sd205   , -10'sd469   }; /* W[ 189] =  0.4004  -0.9160i */
dout[702]= { 10'sd202   , -10'sd471   }; /* W[ 190] =  0.3945  -0.9199i */
dout[703]= { 10'sd199   , -10'sd472   }; /* W[ 191] =  0.3887  -0.9219i */
dout[704]= { 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[705]= { 10'sd193   , -10'sd474   }; /* W[ 193] =  0.3770  -0.9258i */
dout[706]= { 10'sd190   , -10'sd475   }; /* W[ 194] =  0.3711  -0.9277i */
dout[707]= { 10'sd187   , -10'sd477   }; /* W[ 195] =  0.3652  -0.9316i */
dout[708]= { 10'sd184   , -10'sd478   }; /* W[ 196] =  0.3594  -0.9336i */
dout[709]= { 10'sd181   , -10'sd479   }; /* W[ 197] =  0.3535  -0.9355i */
dout[710]= { 10'sd178   , -10'sd480   }; /* W[ 198] =  0.3477  -0.9375i */
dout[711]= { 10'sd175   , -10'sd481   }; /* W[ 199] =  0.3418  -0.9395i */
dout[712]= { 10'sd172   , -10'sd482   }; /* W[ 200] =  0.3359  -0.9414i */
dout[713]= { 10'sd170   , -10'sd483   }; /* W[ 201] =  0.3320  -0.9434i */
dout[714]= { 10'sd167   , -10'sd484   }; /* W[ 202] =  0.3262  -0.9453i */
dout[715]= { 10'sd164   , -10'sd485   }; /* W[ 203] =  0.3203  -0.9473i */
dout[716]= { 10'sd161   , -10'sd486   }; /* W[ 204] =  0.3145  -0.9492i */
dout[717]= { 10'sd158   , -10'sd487   }; /* W[ 205] =  0.3086  -0.9512i */
dout[718]= { 10'sd155   , -10'sd488   }; /* W[ 206] =  0.3027  -0.9531i */
dout[719]= { 10'sd152   , -10'sd489   }; /* W[ 207] =  0.2969  -0.9551i */
dout[720]= { 10'sd149   , -10'sd490   }; /* W[ 208] =  0.2910  -0.9570i */
dout[721]= { 10'sd146   , -10'sd491   }; /* W[ 209] =  0.2852  -0.9590i */
dout[722]= { 10'sd143   , -10'sd492   }; /* W[ 210] =  0.2793  -0.9609i */
dout[723]= { 10'sd140   , -10'sd493   }; /* W[ 211] =  0.2734  -0.9629i */
dout[724]= { 10'sd137   , -10'sd493   }; /* W[ 212] =  0.2676  -0.9629i */
dout[725]= { 10'sd134   , -10'sd494   }; /* W[ 213] =  0.2617  -0.9648i */
dout[726]= { 10'sd130   , -10'sd495   }; /* W[ 214] =  0.2539  -0.9668i */
dout[727]= { 10'sd127   , -10'sd496   }; /* W[ 215] =  0.2480  -0.9688i */
dout[728]= { 10'sd124   , -10'sd497   }; /* W[ 216] =  0.2422  -0.9707i */
dout[729]= { 10'sd121   , -10'sd497   }; /* W[ 217] =  0.2363  -0.9707i */
dout[730]= { 10'sd118   , -10'sd498   }; /* W[ 218] =  0.2305  -0.9727i */
dout[731]= { 10'sd115   , -10'sd499   }; /* W[ 219] =  0.2246  -0.9746i */
dout[732]= { 10'sd112   , -10'sd500   }; /* W[ 220] =  0.2188  -0.9766i */
dout[733]= { 10'sd109   , -10'sd500   }; /* W[ 221] =  0.2129  -0.9766i */
dout[734]= { 10'sd106   , -10'sd501   }; /* W[ 222] =  0.2070  -0.9785i */
dout[735]= { 10'sd103   , -10'sd502   }; /* W[ 223] =  0.2012  -0.9805i */
dout[736]= { 10'sd100   , -10'sd502   }; /* W[ 224] =  0.1953  -0.9805i */
dout[737]= { 10'sd97    , -10'sd503   }; /* W[ 225] =  0.1895  -0.9824i */
dout[738]= { 10'sd94    , -10'sd503   }; /* W[ 226] =  0.1836  -0.9824i */
dout[739]= { 10'sd91    , -10'sd504   }; /* W[ 227] =  0.1777  -0.9844i */
dout[740]= { 10'sd88    , -10'sd504   }; /* W[ 228] =  0.1719  -0.9844i */
dout[741]= { 10'sd84    , -10'sd505   }; /* W[ 229] =  0.1641  -0.9863i */
dout[742]= { 10'sd81    , -10'sd505   }; /* W[ 230] =  0.1582  -0.9863i */
dout[743]= { 10'sd78    , -10'sd506   }; /* W[ 231] =  0.1523  -0.9883i */
dout[744]= { 10'sd75    , -10'sd506   }; /* W[ 232] =  0.1465  -0.9883i */
dout[745]= { 10'sd72    , -10'sd507   }; /* W[ 233] =  0.1406  -0.9902i */
dout[746]= { 10'sd69    , -10'sd507   }; /* W[ 234] =  0.1348  -0.9902i */
dout[747]= { 10'sd66    , -10'sd508   }; /* W[ 235] =  0.1289  -0.9922i */
dout[748]= { 10'sd63    , -10'sd508   }; /* W[ 236] =  0.1230  -0.9922i */
dout[749]= { 10'sd60    , -10'sd509   }; /* W[ 237] =  0.1172  -0.9941i */
dout[750]= { 10'sd56    , -10'sd509   }; /* W[ 238] =  0.1094  -0.9941i */
dout[751]= { 10'sd53    , -10'sd509   }; /* W[ 239] =  0.1035  -0.9941i */
dout[752]= { 10'sd50    , -10'sd510   }; /* W[ 240] =  0.0977  -0.9961i */
dout[753]= { 10'sd47    , -10'sd510   }; /* W[ 241] =  0.0918  -0.9961i */
dout[754]= { 10'sd44    , -10'sd510   }; /* W[ 242] =  0.0859  -0.9961i */
dout[755]= { 10'sd41    , -10'sd510   }; /* W[ 243] =  0.0801  -0.9961i */
dout[756]= { 10'sd38    , -10'sd511   }; /* W[ 244] =  0.0742  -0.9980i */
dout[757]= { 10'sd35    , -10'sd511   }; /* W[ 245] =  0.0684  -0.9980i */
dout[758]= { 10'sd31    , -10'sd511   }; /* W[ 246] =  0.0605  -0.9980i */
dout[759]= { 10'sd28    , -10'sd511   }; /* W[ 247] =  0.0547  -0.9980i */
dout[760]= { 10'sd25    , -10'sd511   }; /* W[ 248] =  0.0488  -0.9980i */
dout[761]= { 10'sd22    , -10'sd512   }; /* W[ 249] =  0.0430  -1.0000i */
dout[762]= { 10'sd19    , -10'sd512   }; /* W[ 250] =  0.0371  -1.0000i */
dout[763]= { 10'sd16    , -10'sd512   }; /* W[ 251] =  0.0312  -1.0000i */
dout[764]= { 10'sd13    , -10'sd512   }; /* W[ 252] =  0.0254  -1.0000i */
dout[765]= { 10'sd9     , -10'sd512   }; /* W[ 253] =  0.0176  -1.0000i */
dout[766]= { 10'sd6     , -10'sd512   }; /* W[ 254] =  0.0117  -1.0000i */
dout[767]= { 10'sd3     , -10'sd512   }; /* W[ 255] =  0.0059  -1.0000i */
dout[768]= { 10'sd511   ,  10'sd0     }; /* W[   0] =  0.9980   0.0000i */
dout[769]= { 10'sd511   , -10'sd9     }; /* W[   3] =  0.9980  -0.0176i */
dout[770]= { 10'sd511   , -10'sd19    }; /* W[   6] =  0.9980  -0.0371i */
dout[771]= { 10'sd511   , -10'sd28    }; /* W[   9] =  0.9980  -0.0547i */
dout[772]= { 10'sd511   , -10'sd38    }; /* W[  12] =  0.9980  -0.0742i */
dout[773]= { 10'sd510   , -10'sd47    }; /* W[  15] =  0.9961  -0.0918i */
dout[774]= { 10'sd509   , -10'sd56    }; /* W[  18] =  0.9941  -0.1094i */
dout[775]= { 10'sd508   , -10'sd66    }; /* W[  21] =  0.9922  -0.1289i */
dout[776]= { 10'sd506   , -10'sd75    }; /* W[  24] =  0.9883  -0.1465i */
dout[777]= { 10'sd505   , -10'sd84    }; /* W[  27] =  0.9863  -0.1641i */
dout[778]= { 10'sd503   , -10'sd94    }; /* W[  30] =  0.9824  -0.1836i */
dout[779]= { 10'sd502   , -10'sd103   }; /* W[  33] =  0.9805  -0.2012i */
dout[780]= { 10'sd500   , -10'sd112   }; /* W[  36] =  0.9766  -0.2188i */
dout[781]= { 10'sd497   , -10'sd121   }; /* W[  39] =  0.9707  -0.2363i */
dout[782]= { 10'sd495   , -10'sd130   }; /* W[  42] =  0.9668  -0.2539i */
dout[783]= { 10'sd493   , -10'sd140   }; /* W[  45] =  0.9629  -0.2734i */
dout[784]= { 10'sd490   , -10'sd149   }; /* W[  48] =  0.9570  -0.2910i */
dout[785]= { 10'sd487   , -10'sd158   }; /* W[  51] =  0.9512  -0.3086i */
dout[786]= { 10'sd484   , -10'sd167   }; /* W[  54] =  0.9453  -0.3262i */
dout[787]= { 10'sd481   , -10'sd175   }; /* W[  57] =  0.9395  -0.3418i */
dout[788]= { 10'sd478   , -10'sd184   }; /* W[  60] =  0.9336  -0.3594i */
dout[789]= { 10'sd474   , -10'sd193   }; /* W[  63] =  0.9258  -0.3770i */
dout[790]= { 10'sd471   , -10'sd202   }; /* W[  66] =  0.9199  -0.3945i */
dout[791]= { 10'sd467   , -10'sd210   }; /* W[  69] =  0.9121  -0.4102i */
dout[792]= { 10'sd463   , -10'sd219   }; /* W[  72] =  0.9043  -0.4277i */
dout[793]= { 10'sd459   , -10'sd227   }; /* W[  75] =  0.8965  -0.4434i */
dout[794]= { 10'sd454   , -10'sd236   }; /* W[  78] =  0.8867  -0.4609i */
dout[795]= { 10'sd450   , -10'sd244   }; /* W[  81] =  0.8789  -0.4766i */
dout[796]= { 10'sd445   , -10'sd252   }; /* W[  84] =  0.8691  -0.4922i */
dout[797]= { 10'sd441   , -10'sd261   }; /* W[  87] =  0.8613  -0.5098i */
dout[798]= { 10'sd436   , -10'sd269   }; /* W[  90] =  0.8516  -0.5254i */
dout[799]= { 10'sd431   , -10'sd277   }; /* W[  93] =  0.8418  -0.5410i */
dout[800]= { 10'sd426   , -10'sd284   }; /* W[  96] =  0.8320  -0.5547i */
dout[801]= { 10'sd420   , -10'sd292   }; /* W[  99] =  0.8203  -0.5703i */
dout[802]= { 10'sd415   , -10'sd300   }; /* W[ 102] =  0.8105  -0.5859i */
dout[803]= { 10'sd409   , -10'sd308   }; /* W[ 105] =  0.7988  -0.6016i */
dout[804]= { 10'sd404   , -10'sd315   }; /* W[ 108] =  0.7891  -0.6152i */
dout[805]= { 10'sd398   , -10'sd322   }; /* W[ 111] =  0.7773  -0.6289i */
dout[806]= { 10'sd392   , -10'sd330   }; /* W[ 114] =  0.7656  -0.6445i */
dout[807]= { 10'sd386   , -10'sd337   }; /* W[ 117] =  0.7539  -0.6582i */
dout[808]= { 10'sd379   , -10'sd344   }; /* W[ 120] =  0.7402  -0.6719i */
dout[809]= { 10'sd373   , -10'sd351   }; /* W[ 123] =  0.7285  -0.6855i */
dout[810]= { 10'sd366   , -10'sd358   }; /* W[ 126] =  0.7148  -0.6992i */
dout[811]= { 10'sd360   , -10'sd364   }; /* W[ 129] =  0.7031  -0.7109i */
dout[812]= { 10'sd353   , -10'sd371   }; /* W[ 132] =  0.6895  -0.7246i */
dout[813]= { 10'sd346   , -10'sd377   }; /* W[ 135] =  0.6758  -0.7363i */
dout[814]= { 10'sd339   , -10'sd384   }; /* W[ 138] =  0.6621  -0.7500i */
dout[815]= { 10'sd332   , -10'sd390   }; /* W[ 141] =  0.6484  -0.7617i */
dout[816]= { 10'sd325   , -10'sd396   }; /* W[ 144] =  0.6348  -0.7734i */
dout[817]= { 10'sd317   , -10'sd402   }; /* W[ 147] =  0.6191  -0.7852i */
dout[818]= { 10'sd310   , -10'sd407   }; /* W[ 150] =  0.6055  -0.7949i */
dout[819]= { 10'sd302   , -10'sd413   }; /* W[ 153] =  0.5898  -0.8066i */
dout[820]= { 10'sd295   , -10'sd419   }; /* W[ 156] =  0.5762  -0.8184i */
dout[821]= { 10'sd287   , -10'sd424   }; /* W[ 159] =  0.5605  -0.8281i */
dout[822]= { 10'sd279   , -10'sd429   }; /* W[ 162] =  0.5449  -0.8379i */
dout[823]= { 10'sd271   , -10'sd434   }; /* W[ 165] =  0.5293  -0.8477i */
dout[824]= { 10'sd263   , -10'sd439   }; /* W[ 168] =  0.5137  -0.8574i */
dout[825]= { 10'sd255   , -10'sd444   }; /* W[ 171] =  0.4980  -0.8672i */
dout[826]= { 10'sd247   , -10'sd449   }; /* W[ 174] =  0.4824  -0.8770i */
dout[827]= { 10'sd239   , -10'sd453   }; /* W[ 177] =  0.4668  -0.8848i */
dout[828]= { 10'sd230   , -10'sd457   }; /* W[ 180] =  0.4492  -0.8926i */
dout[829]= { 10'sd222   , -10'sd461   }; /* W[ 183] =  0.4336  -0.9004i */
dout[830]= { 10'sd213   , -10'sd465   }; /* W[ 186] =  0.4160  -0.9082i */
dout[831]= { 10'sd205   , -10'sd469   }; /* W[ 189] =  0.4004  -0.9160i */
dout[832]= { 10'sd196   , -10'sd473   }; /* W[ 192] =  0.3828  -0.9238i */
dout[833]= { 10'sd187   , -10'sd477   }; /* W[ 195] =  0.3652  -0.9316i */
dout[834]= { 10'sd178   , -10'sd480   }; /* W[ 198] =  0.3477  -0.9375i */
dout[835]= { 10'sd170   , -10'sd483   }; /* W[ 201] =  0.3320  -0.9434i */
dout[836]= { 10'sd161   , -10'sd486   }; /* W[ 204] =  0.3145  -0.9492i */
dout[837]= { 10'sd152   , -10'sd489   }; /* W[ 207] =  0.2969  -0.9551i */
dout[838]= { 10'sd143   , -10'sd492   }; /* W[ 210] =  0.2793  -0.9609i */
dout[839]= { 10'sd134   , -10'sd494   }; /* W[ 213] =  0.2617  -0.9648i */
dout[840]= { 10'sd124   , -10'sd497   }; /* W[ 216] =  0.2422  -0.9707i */
dout[841]= { 10'sd115   , -10'sd499   }; /* W[ 219] =  0.2246  -0.9746i */
dout[842]= { 10'sd106   , -10'sd501   }; /* W[ 222] =  0.2070  -0.9785i */
dout[843]= { 10'sd97    , -10'sd503   }; /* W[ 225] =  0.1895  -0.9824i */
dout[844]= { 10'sd88    , -10'sd504   }; /* W[ 228] =  0.1719  -0.9844i */
dout[845]= { 10'sd78    , -10'sd506   }; /* W[ 231] =  0.1523  -0.9883i */
dout[846]= { 10'sd69    , -10'sd507   }; /* W[ 234] =  0.1348  -0.9902i */
dout[847]= { 10'sd60    , -10'sd509   }; /* W[ 237] =  0.1172  -0.9941i */
dout[848]= { 10'sd50    , -10'sd510   }; /* W[ 240] =  0.0977  -0.9961i */
dout[849]= { 10'sd41    , -10'sd510   }; /* W[ 243] =  0.0801  -0.9961i */
dout[850]= { 10'sd31    , -10'sd511   }; /* W[ 246] =  0.0605  -0.9980i */
dout[851]= { 10'sd22    , -10'sd512   }; /* W[ 249] =  0.0430  -1.0000i */
dout[852]= { 10'sd13    , -10'sd512   }; /* W[ 252] =  0.0254  -1.0000i */
dout[853]= { 10'sd3     , -10'sd512   }; /* W[ 255] =  0.0059  -1.0000i */
dout[854]= {-10'sd6     , -10'sd512   }; /* W[ 258] = -0.0117  -1.0000i */
dout[855]= {-10'sd16    , -10'sd512   }; /* W[ 261] = -0.0312  -1.0000i */
dout[856]= {-10'sd25    , -10'sd511   }; /* W[ 264] = -0.0488  -0.9980i */
dout[857]= {-10'sd35    , -10'sd511   }; /* W[ 267] = -0.0684  -0.9980i */
dout[858]= {-10'sd44    , -10'sd510   }; /* W[ 270] = -0.0859  -0.9961i */
dout[859]= {-10'sd53    , -10'sd509   }; /* W[ 273] = -0.1035  -0.9941i */
dout[860]= {-10'sd63    , -10'sd508   }; /* W[ 276] = -0.1230  -0.9922i */
dout[861]= {-10'sd72    , -10'sd507   }; /* W[ 279] = -0.1406  -0.9902i */
dout[862]= {-10'sd81    , -10'sd505   }; /* W[ 282] = -0.1582  -0.9863i */
dout[863]= {-10'sd91    , -10'sd504   }; /* W[ 285] = -0.1777  -0.9844i */
dout[864]= {-10'sd100   , -10'sd502   }; /* W[ 288] = -0.1953  -0.9805i */
dout[865]= {-10'sd109   , -10'sd500   }; /* W[ 291] = -0.2129  -0.9766i */
dout[866]= {-10'sd118   , -10'sd498   }; /* W[ 294] = -0.2305  -0.9727i */
dout[867]= {-10'sd127   , -10'sd496   }; /* W[ 297] = -0.2480  -0.9688i */
dout[868]= {-10'sd137   , -10'sd493   }; /* W[ 300] = -0.2676  -0.9629i */
dout[869]= {-10'sd146   , -10'sd491   }; /* W[ 303] = -0.2852  -0.9590i */
dout[870]= {-10'sd155   , -10'sd488   }; /* W[ 306] = -0.3027  -0.9531i */
dout[871]= {-10'sd164   , -10'sd485   }; /* W[ 309] = -0.3203  -0.9473i */
dout[872]= {-10'sd172   , -10'sd482   }; /* W[ 312] = -0.3359  -0.9414i */
dout[873]= {-10'sd181   , -10'sd479   }; /* W[ 315] = -0.3535  -0.9355i */
dout[874]= {-10'sd190   , -10'sd475   }; /* W[ 318] = -0.3711  -0.9277i */
dout[875]= {-10'sd199   , -10'sd472   }; /* W[ 321] = -0.3887  -0.9219i */
dout[876]= {-10'sd207   , -10'sd468   }; /* W[ 324] = -0.4043  -0.9141i */
dout[877]= {-10'sd216   , -10'sd464   }; /* W[ 327] = -0.4219  -0.9062i */
dout[878]= {-10'sd225   , -10'sd460   }; /* W[ 330] = -0.4395  -0.8984i */
dout[879]= {-10'sd233   , -10'sd456   }; /* W[ 333] = -0.4551  -0.8906i */
dout[880]= {-10'sd241   , -10'sd452   }; /* W[ 336] = -0.4707  -0.8828i */
dout[881]= {-10'sd250   , -10'sd447   }; /* W[ 339] = -0.4883  -0.8730i */
dout[882]= {-10'sd258   , -10'sd442   }; /* W[ 342] = -0.5039  -0.8633i */
dout[883]= {-10'sd266   , -10'sd438   }; /* W[ 345] = -0.5195  -0.8555i */
dout[884]= {-10'sd274   , -10'sd433   }; /* W[ 348] = -0.5352  -0.8457i */
dout[885]= {-10'sd282   , -10'sd427   }; /* W[ 351] = -0.5508  -0.8340i */
dout[886]= {-10'sd290   , -10'sd422   }; /* W[ 354] = -0.5664  -0.8242i */
dout[887]= {-10'sd297   , -10'sd417   }; /* W[ 357] = -0.5801  -0.8145i */
dout[888]= {-10'sd305   , -10'sd411   }; /* W[ 360] = -0.5957  -0.8027i */
dout[889]= {-10'sd313   , -10'sd406   }; /* W[ 363] = -0.6113  -0.7930i */
dout[890]= {-10'sd320   , -10'sd400   }; /* W[ 366] = -0.6250  -0.7812i */
dout[891]= {-10'sd327   , -10'sd394   }; /* W[ 369] = -0.6387  -0.7695i */
dout[892]= {-10'sd334   , -10'sd388   }; /* W[ 372] = -0.6523  -0.7578i */
dout[893]= {-10'sd342   , -10'sd381   }; /* W[ 375] = -0.6680  -0.7441i */
dout[894]= {-10'sd348   , -10'sd375   }; /* W[ 378] = -0.6797  -0.7324i */
dout[895]= {-10'sd355   , -10'sd369   }; /* W[ 381] = -0.6934  -0.7207i */
dout[896]= {-10'sd362   , -10'sd362   }; /* W[ 384] = -0.7070  -0.7070i */
dout[897]= {-10'sd369   , -10'sd355   }; /* W[ 387] = -0.7207  -0.6934i */
dout[898]= {-10'sd375   , -10'sd348   }; /* W[ 390] = -0.7324  -0.6797i */
dout[899]= {-10'sd381   , -10'sd342   }; /* W[ 393] = -0.7441  -0.6680i */
dout[900]= {-10'sd388   , -10'sd334   }; /* W[ 396] = -0.7578  -0.6523i */
dout[901]= {-10'sd394   , -10'sd327   }; /* W[ 399] = -0.7695  -0.6387i */
dout[902]= {-10'sd400   , -10'sd320   }; /* W[ 402] = -0.7812  -0.6250i */
dout[903]= {-10'sd406   , -10'sd313   }; /* W[ 405] = -0.7930  -0.6113i */
dout[904]= {-10'sd411   , -10'sd305   }; /* W[ 408] = -0.8027  -0.5957i */
dout[905]= {-10'sd417   , -10'sd297   }; /* W[ 411] = -0.8145  -0.5801i */
dout[906]= {-10'sd422   , -10'sd290   }; /* W[ 414] = -0.8242  -0.5664i */
dout[907]= {-10'sd427   , -10'sd282   }; /* W[ 417] = -0.8340  -0.5508i */
dout[908]= {-10'sd433   , -10'sd274   }; /* W[ 420] = -0.8457  -0.5352i */
dout[909]= {-10'sd438   , -10'sd266   }; /* W[ 423] = -0.8555  -0.5195i */
dout[910]= {-10'sd442   , -10'sd258   }; /* W[ 426] = -0.8633  -0.5039i */
dout[911]= {-10'sd447   , -10'sd250   }; /* W[ 429] = -0.8730  -0.4883i */
dout[912]= {-10'sd452   , -10'sd241   }; /* W[ 432] = -0.8828  -0.4707i */
dout[913]= {-10'sd456   , -10'sd233   }; /* W[ 435] = -0.8906  -0.4551i */
dout[914]= {-10'sd460   , -10'sd225   }; /* W[ 438] = -0.8984  -0.4395i */
dout[915]= {-10'sd464   , -10'sd216   }; /* W[ 441] = -0.9062  -0.4219i */
dout[916]= {-10'sd468   , -10'sd207   }; /* W[ 444] = -0.9141  -0.4043i */
dout[917]= {-10'sd472   , -10'sd199   }; /* W[ 447] = -0.9219  -0.3887i */
dout[918]= {-10'sd475   , -10'sd190   }; /* W[ 450] = -0.9277  -0.3711i */
dout[919]= {-10'sd479   , -10'sd181   }; /* W[ 453] = -0.9355  -0.3535i */
dout[920]= {-10'sd482   , -10'sd172   }; /* W[ 456] = -0.9414  -0.3359i */
dout[921]= {-10'sd485   , -10'sd164   }; /* W[ 459] = -0.9473  -0.3203i */
dout[922]= {-10'sd488   , -10'sd155   }; /* W[ 462] = -0.9531  -0.3027i */
dout[923]= {-10'sd491   , -10'sd146   }; /* W[ 465] = -0.9590  -0.2852i */
dout[924]= {-10'sd493   , -10'sd137   }; /* W[ 468] = -0.9629  -0.2676i */
dout[925]= {-10'sd496   , -10'sd127   }; /* W[ 471] = -0.9688  -0.2480i */
dout[926]= {-10'sd498   , -10'sd118   }; /* W[ 474] = -0.9727  -0.2305i */
dout[927]= {-10'sd500   , -10'sd109   }; /* W[ 477] = -0.9766  -0.2129i */
dout[928]= {-10'sd502   , -10'sd100   }; /* W[ 480] = -0.9805  -0.1953i */
dout[929]= {-10'sd504   , -10'sd91    }; /* W[ 483] = -0.9844  -0.1777i */
dout[930]= {-10'sd505   , -10'sd81    }; /* W[ 486] = -0.9863  -0.1582i */
dout[931]= {-10'sd507   , -10'sd72    }; /* W[ 489] = -0.9902  -0.1406i */
dout[932]= {-10'sd508   , -10'sd63    }; /* W[ 492] = -0.9922  -0.1230i */
dout[933]= {-10'sd509   , -10'sd53    }; /* W[ 495] = -0.9941  -0.1035i */
dout[934]= {-10'sd510   , -10'sd44    }; /* W[ 498] = -0.9961  -0.0859i */
dout[935]= {-10'sd511   , -10'sd35    }; /* W[ 501] = -0.9980  -0.0684i */
dout[936]= {-10'sd511   , -10'sd25    }; /* W[ 504] = -0.9980  -0.0488i */
dout[937]= {-10'sd512   , -10'sd16    }; /* W[ 507] = -1.0000  -0.0312i */
dout[938]= {-10'sd512   , -10'sd6     }; /* W[ 510] = -1.0000  -0.0117i */
dout[939]= {-10'sd512   ,  10'sd3     }; /* W[ 513] = -1.0000   0.0059i */
dout[940]= {-10'sd512   ,  10'sd13    }; /* W[ 516] = -1.0000   0.0254i */
dout[941]= {-10'sd512   ,  10'sd22    }; /* W[ 519] = -1.0000   0.0430i */
dout[942]= {-10'sd511   ,  10'sd31    }; /* W[ 522] = -0.9980   0.0605i */
dout[943]= {-10'sd510   ,  10'sd41    }; /* W[ 525] = -0.9961   0.0801i */
dout[944]= {-10'sd510   ,  10'sd50    }; /* W[ 528] = -0.9961   0.0977i */
dout[945]= {-10'sd509   ,  10'sd60    }; /* W[ 531] = -0.9941   0.1172i */
dout[946]= {-10'sd507   ,  10'sd69    }; /* W[ 534] = -0.9902   0.1348i */
dout[947]= {-10'sd506   ,  10'sd78    }; /* W[ 537] = -0.9883   0.1523i */
dout[948]= {-10'sd504   ,  10'sd88    }; /* W[ 540] = -0.9844   0.1719i */
dout[949]= {-10'sd503   ,  10'sd97    }; /* W[ 543] = -0.9824   0.1895i */
dout[950]= {-10'sd501   ,  10'sd106   }; /* W[ 546] = -0.9785   0.2070i */
dout[951]= {-10'sd499   ,  10'sd115   }; /* W[ 549] = -0.9746   0.2246i */
dout[952]= {-10'sd497   ,  10'sd124   }; /* W[ 552] = -0.9707   0.2422i */
dout[953]= {-10'sd494   ,  10'sd134   }; /* W[ 555] = -0.9648   0.2617i */
dout[954]= {-10'sd492   ,  10'sd143   }; /* W[ 558] = -0.9609   0.2793i */
dout[955]= {-10'sd489   ,  10'sd152   }; /* W[ 561] = -0.9551   0.2969i */
dout[956]= {-10'sd486   ,  10'sd161   }; /* W[ 564] = -0.9492   0.3145i */
dout[957]= {-10'sd483   ,  10'sd170   }; /* W[ 567] = -0.9434   0.3320i */
dout[958]= {-10'sd480   ,  10'sd178   }; /* W[ 570] = -0.9375   0.3477i */
dout[959]= {-10'sd477   ,  10'sd187   }; /* W[ 573] = -0.9316   0.3652i */
dout[960]= {-10'sd473   ,  10'sd196   }; /* W[ 576] = -0.9238   0.3828i */
dout[961]= {-10'sd469   ,  10'sd205   }; /* W[ 579] = -0.9160   0.4004i */
dout[962]= {-10'sd465   ,  10'sd213   }; /* W[ 582] = -0.9082   0.4160i */
dout[963]= {-10'sd461   ,  10'sd222   }; /* W[ 585] = -0.9004   0.4336i */
dout[964]= {-10'sd457   ,  10'sd230   }; /* W[ 588] = -0.8926   0.4492i */
dout[965]= {-10'sd453   ,  10'sd239   }; /* W[ 591] = -0.8848   0.4668i */
dout[966]= {-10'sd449   ,  10'sd247   }; /* W[ 594] = -0.8770   0.4824i */
dout[967]= {-10'sd444   ,  10'sd255   }; /* W[ 597] = -0.8672   0.4980i */
dout[968]= {-10'sd439   ,  10'sd263   }; /* W[ 600] = -0.8574   0.5137i */
dout[969]= {-10'sd434   ,  10'sd271   }; /* W[ 603] = -0.8477   0.5293i */
dout[970]= {-10'sd429   ,  10'sd279   }; /* W[ 606] = -0.8379   0.5449i */
dout[971]= {-10'sd424   ,  10'sd287   }; /* W[ 609] = -0.8281   0.5605i */
dout[972]= {-10'sd419   ,  10'sd295   }; /* W[ 612] = -0.8184   0.5762i */
dout[973]= {-10'sd413   ,  10'sd302   }; /* W[ 615] = -0.8066   0.5898i */
dout[974]= {-10'sd407   ,  10'sd310   }; /* W[ 618] = -0.7949   0.6055i */
dout[975]= {-10'sd402   ,  10'sd317   }; /* W[ 621] = -0.7852   0.6191i */
dout[976]= {-10'sd396   ,  10'sd325   }; /* W[ 624] = -0.7734   0.6348i */
dout[977]= {-10'sd390   ,  10'sd332   }; /* W[ 627] = -0.7617   0.6484i */
dout[978]= {-10'sd384   ,  10'sd339   }; /* W[ 630] = -0.7500   0.6621i */
dout[979]= {-10'sd377   ,  10'sd346   }; /* W[ 633] = -0.7363   0.6758i */
dout[980]= {-10'sd371   ,  10'sd353   }; /* W[ 636] = -0.7246   0.6895i */
dout[981]= {-10'sd364   ,  10'sd360   }; /* W[ 639] = -0.7109   0.7031i */
dout[982]= {-10'sd358   ,  10'sd366   }; /* W[ 642] = -0.6992   0.7148i */
dout[983]= {-10'sd351   ,  10'sd373   }; /* W[ 645] = -0.6855   0.7285i */
dout[984]= {-10'sd344   ,  10'sd379   }; /* W[ 648] = -0.6719   0.7402i */
dout[985]= {-10'sd337   ,  10'sd386   }; /* W[ 651] = -0.6582   0.7539i */
dout[986]= {-10'sd330   ,  10'sd392   }; /* W[ 654] = -0.6445   0.7656i */
dout[987]= {-10'sd322   ,  10'sd398   }; /* W[ 657] = -0.6289   0.7773i */
dout[988]= {-10'sd315   ,  10'sd404   }; /* W[ 660] = -0.6152   0.7891i */
dout[989]= {-10'sd308   ,  10'sd409   }; /* W[ 663] = -0.6016   0.7988i */
dout[990]= {-10'sd300   ,  10'sd415   }; /* W[ 666] = -0.5859   0.8105i */
dout[991]= {-10'sd292   ,  10'sd420   }; /* W[ 669] = -0.5703   0.8203i */
dout[992]= {-10'sd284   ,  10'sd426   }; /* W[ 672] = -0.5547   0.8320i */
dout[993]= {-10'sd277   ,  10'sd431   }; /* W[ 675] = -0.5410   0.8418i */
dout[994]= {-10'sd269   ,  10'sd436   }; /* W[ 678] = -0.5254   0.8516i */
dout[995]= {-10'sd261   ,  10'sd441   }; /* W[ 681] = -0.5098   0.8613i */
dout[996]= {-10'sd252   ,  10'sd445   }; /* W[ 684] = -0.4922   0.8691i */
dout[997]= {-10'sd244   ,  10'sd450   }; /* W[ 687] = -0.4766   0.8789i */
dout[998]= {-10'sd236   ,  10'sd454   }; /* W[ 690] = -0.4609   0.8867i */
dout[999]= {-10'sd227   ,  10'sd459   }; /* W[ 693] = -0.4434   0.8965i */
dout[1000]= {-10'sd219   ,  10'sd463   }; /* W[ 696] = -0.4277   0.9043i */
dout[1001]= {-10'sd210   ,  10'sd467   }; /* W[ 699] = -0.4102   0.9121i */
dout[1002]= {-10'sd202   ,  10'sd471   }; /* W[ 702] = -0.3945   0.9199i */
dout[1003]= {-10'sd193   ,  10'sd474   }; /* W[ 705] = -0.3770   0.9258i */
dout[1004]= {-10'sd184   ,  10'sd478   }; /* W[ 708] = -0.3594   0.9336i */
dout[1005]= {-10'sd175   ,  10'sd481   }; /* W[ 711] = -0.3418   0.9395i */
dout[1006]= {-10'sd167   ,  10'sd484   }; /* W[ 714] = -0.3262   0.9453i */
dout[1007]= {-10'sd158   ,  10'sd487   }; /* W[ 717] = -0.3086   0.9512i */
dout[1008]= {-10'sd149   ,  10'sd490   }; /* W[ 720] = -0.2910   0.9570i */
dout[1009]= {-10'sd140   ,  10'sd493   }; /* W[ 723] = -0.2734   0.9629i */
dout[1010]= {-10'sd130   ,  10'sd495   }; /* W[ 726] = -0.2539   0.9668i */
dout[1011]= {-10'sd121   ,  10'sd497   }; /* W[ 729] = -0.2363   0.9707i */
dout[1012]= {-10'sd112   ,  10'sd500   }; /* W[ 732] = -0.2188   0.9766i */
dout[1013]= {-10'sd103   ,  10'sd502   }; /* W[ 735] = -0.2012   0.9805i */
dout[1014]= {-10'sd94    ,  10'sd503   }; /* W[ 738] = -0.1836   0.9824i */
dout[1015]= {-10'sd84    ,  10'sd505   }; /* W[ 741] = -0.1641   0.9863i */
dout[1016]= {-10'sd75    ,  10'sd506   }; /* W[ 744] = -0.1465   0.9883i */
dout[1017]= {-10'sd66    ,  10'sd508   }; /* W[ 747] = -0.1289   0.9922i */
dout[1018]= {-10'sd56    ,  10'sd509   }; /* W[ 750] = -0.1094   0.9941i */
dout[1019]= {-10'sd47    ,  10'sd510   }; /* W[ 753] = -0.0918   0.9961i */
dout[1020]= {-10'sd38    ,  10'sd511   }; /* W[ 756] = -0.0742   0.9980i */
dout[1021]= {-10'sd28    ,  10'sd511   }; /* W[ 759] = -0.0547   0.9980i */
dout[1022]= {-10'sd19    ,  10'sd511   }; /* W[ 762] = -0.0371   0.9980i */
dout[1023]= {-10'sd9     ,  10'sd511   }; /* W[ 765] = -0.0176   0.9980i */
end

always @ (posedge clk) begin
  tf_re<=dout[addr][19:10];
  tf_im<=dout[addr][9:0];
end


endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */
