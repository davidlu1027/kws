module kernel_3_rom (
    input  wire        [ 7:0] addr,
    input  wire               in_valid,
    input  wire               clk,
    output reg signed [ 191:0] w
  );

reg [191:0] dout [0:143];


initial begin
dout[0]={ -16'd8525,16'd10654,16'd3928,-16'd6242,-16'd13794,-16'd9925,-16'd9891,16'd3101,-16'd8647,-16'd5221,16'd8203,-16'd7607};
dout[1]={ 16'd6808,16'd2516,16'd1159,16'd3161,16'd3012,16'd159,16'd10119,16'd7845,-16'd4714,-16'd2824,16'd11758,16'd9184};
dout[2]={ -16'd3485,-16'd8562,16'd8131,-16'd6853,-16'd1644,16'd10877,16'd7018,-16'd3023,16'd12198,-16'd11372,-16'd3234,16'd9345};
dout[3]={ -16'd1775,-16'd5507,16'd4791,-16'd6853,-16'd2235,-16'd445,16'd1203,16'd5170,-16'd10818,-16'd10047,16'd9048,-16'd1394};
dout[4]={ -16'd12520,16'd8206,-16'd9334,-16'd8318,-16'd2514,-16'd7770,-16'd3270,-16'd5733,16'd6472,16'd7584,-16'd1369,-16'd4696};
dout[5]={ -16'd15269,16'd1742,16'd9019,16'd9506,16'd544,16'd10370,-16'd8300,-16'd10725,-16'd10363,-16'd9446,16'd537,-16'd433};
dout[6]={ 16'd8505,16'd4786,16'd6930,16'd8656,16'd1718,16'd11869,16'd5709,16'd3722,16'd4318,16'd2889,-16'd2225,16'd3427};
dout[7]={ -16'd6791,16'd4652,16'd4715,-16'd11206,16'd9105,-16'd11639,16'd10485,-16'd2293,16'd4657,-16'd7712,-16'd5877,16'd5976};
dout[8]={ -16'd3405,16'd11984,-16'd7941,-16'd5388,-16'd8049,-16'd4375,16'd4932,16'd11960,-16'd5792,-16'd4870,16'd2305,-16'd7189};
dout[9]={ 16'd15264,16'd8340,16'd1481,-16'd1711,16'd6629,-16'd10445,-16'd3557,-16'd10417,16'd1415,16'd2252,-16'd251,16'd4116};
dout[10]={ -16'd4532,-16'd8337,16'd10975,-16'd11535,16'd1394,16'd8113,-16'd12611,16'd1172,16'd5856,-16'd7086,-16'd2813,16'd8124};
dout[11]={ 16'd41953,-16'd11809,-16'd11666,-16'd5373,16'd7254,-16'd7374,-16'd10318,-16'd11601,16'd9119,16'd7521,16'd4278,-16'd22672};
dout[12]={ 16'd35090,-16'd7507,-16'd5397,-16'd14704,-16'd631,16'd3450,-16'd13043,-16'd1521,-16'd18856,-16'd12108,-16'd2434,-16'd13897};
dout[13]={ -16'd25006,16'd9839,16'd55,-16'd11799,-16'd6116,-16'd9671,16'd3591,-16'd725,-16'd993,-16'd7748,16'd3176,-16'd4713};
dout[14]={ -16'd16366,16'd5584,-16'd13601,16'd10563,-16'd3319,16'd12887,-16'd10723,-16'd2535,-16'd9714,-16'd6530,16'd11382,16'd3833};
dout[15]={ -16'd5706,-16'd3682,-16'd4939,-16'd2736,-16'd7075,16'd5751,-16'd4589,16'd3837,-16'd5252,-16'd6134,-16'd7913,16'd7767};
dout[16]={ -16'd6664,-16'd5266,-16'd895,-16'd7205,16'd11408,-16'd9098,16'd2926,-16'd8397,16'd6008,-16'd8623,-16'd12452,-16'd7106};
dout[17]={ -16'd14616,-16'd1079,-16'd5021,16'd4210,-16'd3832,16'd5310,16'd727,-16'd8587,-16'd6585,16'd562,-16'd2309,16'd1642};
dout[18]={ 16'd8613,-16'd7777,16'd2788,-16'd7054,16'd7419,-16'd2626,16'd2171,-16'd9607,-16'd9459,-16'd7766,-16'd7288,16'd3120};
dout[19]={ -16'd498,16'd11756,-16'd6175,16'd1709,-16'd4524,-16'd8319,16'd9934,-16'd1869,16'd6966,16'd5947,16'd5010,16'd8206};
dout[20]={ 16'd4663,-16'd8113,16'd7523,16'd3519,-16'd5461,-16'd4724,16'd4798,16'd2307,-16'd11758,16'd9460,16'd10645,16'd4357};
dout[21]={ 16'd2171,16'd5595,16'd10262,16'd2742,16'd5003,-16'd2086,16'd8722,16'd13785,16'd4354,16'd3267,-16'd2401,-16'd5703};
dout[22]={ -16'd22587,-16'd2663,16'd4998,-16'd1841,-16'd15358,16'd7517,-16'd14077,16'd3412,-16'd2196,-16'd5065,16'd2888,16'd3806};
dout[23]={ 16'd4719,-16'd1464,-16'd7944,-16'd2266,16'd2706,-16'd367,-16'd10213,-16'd7136,16'd3846,16'd8498,-16'd4817,-16'd3050};
dout[24]={ 16'd15910,-16'd2779,-16'd338,16'd7331,16'd4292,-16'd4242,-16'd9075,-16'd9851,-16'd12095,-16'd2299,16'd288,16'd7122};
dout[25]={ -16'd3374,-16'd6957,-16'd5636,16'd9512,-16'd9739,-16'd7276,-16'd950,-16'd6622,-16'd12288,16'd6368,16'd12272,-16'd406};
dout[26]={ -16'd11393,16'd236,-16'd4154,-16'd8554,-16'd694,-16'd9322,16'd3334,16'd12758,16'd2190,-16'd1393,16'd4853,-16'd6041};
dout[27]={ -16'd9563,16'd10634,16'd2774,16'd8700,16'd6524,16'd3622,16'd11740,16'd6602,16'd3815,16'd12340,16'd10891,16'd9638};
dout[28]={ -16'd4946,16'd2807,-16'd4717,16'd3370,16'd6876,16'd5213,-16'd6167,16'd7223,16'd9465,-16'd4005,-16'd205,16'd11437};
dout[29]={ 16'd8087,16'd1409,-16'd9824,-16'd6035,16'd8559,-16'd7363,-16'd1901,-16'd964,-16'd7539,-16'd7675,-16'd8762,-16'd8013};
dout[30]={ -16'd14912,-16'd29,16'd5388,-16'd3146,-16'd4956,16'd4513,16'd4126,-16'd7159,-16'd11180,-16'd795,16'd4976,16'd234};
dout[31]={ 16'd6708,-16'd1812,-16'd1938,16'd2761,-16'd3225,-16'd3316,-16'd4846,16'd5574,-16'd543,-16'd9045,-16'd1268,16'd5285};
dout[32]={ -16'd7033,16'd9540,16'd3487,16'd3,-16'd6351,-16'd8263,16'd1766,-16'd10161,-16'd6613,-16'd2481,16'd10789,16'd7490};
dout[33]={ 16'd15672,-16'd1187,-16'd10437,16'd5171,-16'd2282,16'd8652,16'd4829,-16'd149,16'd5737,-16'd6614,-16'd5618,16'd6791};
dout[34]={ 16'd14742,16'd7255,16'd8812,-16'd3684,16'd8841,-16'd4717,16'd361,16'd9769,16'd4124,16'd4545,16'd10876,16'd7554};
dout[35]={ 16'd28918,-16'd6260,16'd4538,-16'd770,-16'd2846,-16'd8351,-16'd414,-16'd5198,-16'd8458,-16'd5740,-16'd5365,-16'd5026};
dout[36]={ 16'd7549,16'd2922,16'd5485,-16'd3708,16'd9510,16'd9814,16'd8788,-16'd8029,-16'd3544,-16'd8252,-16'd8701,-16'd2531};
dout[37]={ -16'd8906,-16'd2206,16'd5550,16'd2038,-16'd2504,16'd8210,16'd4666,16'd3820,-16'd1776,-16'd4895,-16'd4969,-16'd6297};
dout[38]={ -16'd10134,16'd2706,16'd10736,16'd8562,16'd850,-16'd645,16'd7505,-16'd10026,16'd5772,-16'd7795,16'd2571,16'd2661};
dout[39]={ -16'd6761,-16'd7734,16'd7962,-16'd1717,-16'd9542,16'd10176,-16'd5677,-16'd13022,-16'd11452,16'd4079,-16'd3144,-16'd2698};
dout[40]={ 16'd10343,-16'd7015,-16'd11383,-16'd724,-16'd2939,-16'd9778,-16'd7051,16'd1362,-16'd10048,-16'd5673,16'd9456,-16'd5994};
dout[41]={ -16'd1662,16'd2733,-16'd7521,-16'd2242,-16'd7247,-16'd9687,16'd4594,16'd5216,16'd67,16'd7993,-16'd1163,-16'd2411};
dout[42]={ -16'd9895,16'd3527,-16'd14976,-16'd10584,16'd1441,-16'd5657,-16'd8075,-16'd6031,-16'd11802,-16'd31,-16'd3838,-16'd5262};
dout[43]={ 16'd12893,16'd710,16'd1978,16'd3918,16'd12556,-16'd12365,-16'd6247,-16'd7502,-16'd3925,16'd4165,16'd6668,16'd2604};
dout[44]={ 16'd28226,16'd4865,-16'd13146,-16'd14483,-16'd13983,-16'd9115,-16'd2027,16'd1053,16'd2742,-16'd9431,16'd6184,-16'd10133};
dout[45]={ -16'd11220,16'd3439,-16'd453,-16'd5962,16'd5811,-16'd6073,16'd3405,16'd3543,-16'd8776,-16'd499,-16'd2729,-16'd5862};
dout[46]={ 16'd7521,-16'd8681,-16'd3702,16'd10081,16'd848,-16'd2324,16'd1001,-16'd11485,-16'd11915,-16'd5283,16'd3167,16'd2761};
dout[47]={ 16'd4377,-16'd4566,16'd15027,16'd9559,16'd11885,-16'd9959,16'd12754,16'd4422,16'd6526,16'd9397,16'd9189,16'd50};
dout[48]={ -16'd3509,16'd427,16'd3875,-16'd9862,16'd7512,-16'd9871,-16'd7962,-16'd11529,16'd9786,16'd9458,-16'd1471,16'd4297};
dout[49]={ -16'd9304,16'd464,-16'd4193,-16'd4772,-16'd7670,16'd1171,16'd5402,16'd2402,16'd11638,-16'd2287,16'd9656,16'd5150};
dout[50]={ 16'd2799,16'd3238,16'd5323,-16'd2664,-16'd4129,16'd689,-16'd132,-16'd1918,16'd8800,16'd13258,-16'd7375,-16'd4482};
dout[51]={ -16'd329,16'd9657,-16'd8761,-16'd4329,16'd8069,-16'd3215,16'd5186,16'd560,16'd2899,-16'd6911,16'd6688,-16'd1691};
dout[52]={ -16'd13970,16'd5048,16'd6349,16'd6532,-16'd4460,16'd949,-16'd1508,16'd350,-16'd10526,-16'd8421,16'd6220,16'd7646};
dout[53]={ -16'd12328,16'd834,16'd296,16'd6508,16'd7368,-16'd47,16'd6696,16'd11311,16'd12092,16'd10949,-16'd4194,16'd12174};
dout[54]={ 16'd15105,16'd5058,16'd2036,16'd4975,16'd4124,16'd3604,16'd9118,-16'd6965,-16'd4751,-16'd10317,-16'd2740,-16'd4171};
dout[55]={ -16'd11211,16'd4212,-16'd8968,16'd4907,-16'd3602,16'd9990,16'd780,16'd3605,-16'd3332,-16'd11186,-16'd2125,-16'd2407};
dout[56]={ 16'd19536,-16'd11346,-16'd2391,16'd3709,-16'd2418,16'd5630,16'd11817,16'd2922,-16'd7736,16'd8703,-16'd10778,-16'd5651};
dout[57]={ -16'd6344,-16'd1142,16'd8598,-16'd5712,16'd4273,-16'd11348,16'd8639,16'd5023,-16'd839,16'd5327,-16'd1878,-16'd9462};
dout[58]={ -16'd4357,16'd8600,16'd3774,-16'd2778,16'd11512,16'd3859,16'd7460,-16'd3929,16'd2303,-16'd1522,-16'd10158,16'd6523};
dout[59]={ -16'd2194,16'd6186,16'd5420,16'd5889,16'd10348,-16'd11357,16'd1363,16'd8895,16'd754,-16'd11074,-16'd8960,16'd4443};
dout[60]={ -16'd20739,-16'd1025,-16'd5891,16'd12031,16'd8049,16'd250,-16'd1880,-16'd3045,-16'd153,-16'd6022,-16'd6764,16'd6204};
dout[61]={ -16'd2883,16'd11136,16'd2971,-16'd1795,16'd8877,16'd2497,-16'd4807,-16'd972,16'd10048,16'd5147,16'd12363,16'd3456};
dout[62]={ -16'd4299,16'd4018,16'd6238,16'd1850,-16'd6843,16'd2670,-16'd6398,-16'd8160,-16'd3070,-16'd9451,16'd8,16'd8691};
dout[63]={ 16'd6187,16'd1752,16'd6132,-16'd3505,-16'd7536,-16'd2319,-16'd1013,16'd8693,-16'd4435,-16'd3265,16'd6993,16'd875};
dout[64]={ -16'd9733,-16'd4225,-16'd1087,16'd3734,16'd4497,16'd6343,16'd1604,-16'd10115,-16'd10331,16'd6718,16'd3014,16'd6932};
dout[65]={ 16'd16153,-16'd4546,16'd2783,-16'd5980,16'd7420,16'd8230,-16'd2551,16'd1089,16'd1496,-16'd5372,16'd8822,16'd5257};
dout[66]={ 16'd6817,16'd5608,16'd896,16'd5333,-16'd6505,16'd3951,-16'd1336,-16'd5331,16'd611,16'd7125,-16'd8386,16'd1852};
dout[67]={ -16'd10111,-16'd4506,-16'd9397,16'd1437,-16'd6258,16'd887,16'd10157,16'd6127,-16'd5059,16'd1931,16'd10501,16'd2211};
dout[68]={ 16'd16844,16'd6689,16'd11075,-16'd11209,-16'd3416,-16'd10112,16'd11865,-16'd8206,-16'd3760,16'd8426,-16'd9003,16'd10772};
dout[69]={ 16'd23172,16'd9887,-16'd15470,-16'd5258,-16'd4306,16'd9646,-16'd11760,-16'd5648,16'd9267,16'd6094,16'd1323,-16'd4590};
dout[70]={ 16'd14694,16'd8625,16'd8128,-16'd5591,16'd3475,-16'd7931,16'd5054,16'd13433,-16'd9997,-16'd7028,-16'd2001,-16'd5669};
dout[71]={ 16'd17585,16'd3956,16'd461,16'd10813,-16'd10543,-16'd7753,-16'd7465,16'd2562,-16'd11127,-16'd11182,-16'd10473,16'd2143};
dout[72]={ 16'd8012,-16'd1667,-16'd8832,-16'd731,16'd9412,16'd6562,16'd5501,-16'd11719,16'd13163,16'd6964,16'd3647,-16'd4246};
dout[73]={ -16'd17000,-16'd6840,-16'd4348,16'd9327,-16'd5883,16'd8293,-16'd8637,-16'd5719,16'd588,16'd2253,-16'd7100,16'd8227};
dout[74]={ -16'd9655,-16'd9599,16'd7081,16'd6880,-16'd7928,-16'd9752,-16'd10690,16'd12250,16'd12437,-16'd6885,-16'd5604,-16'd6311};
dout[75]={ 16'd9816,-16'd7452,-16'd2917,16'd3352,-16'd4233,16'd5367,-16'd1909,-16'd10204,-16'd4122,-16'd7859,-16'd4935,16'd5592};
dout[76]={ -16'd6805,-16'd7953,-16'd2222,-16'd6812,16'd2686,16'd9735,-16'd8356,-16'd5798,-16'd1779,16'd3567,-16'd3054,16'd8148};
dout[77]={ -16'd19060,16'd7290,16'd2559,-16'd1950,16'd3946,-16'd7619,-16'd9842,16'd3881,16'd15846,16'd8677,16'd8698,16'd6370};
dout[78]={ 16'd6500,16'd2446,16'd2728,-16'd12027,-16'd12873,16'd1553,16'd880,16'd6722,16'd3802,-16'd9849,-16'd6370,-16'd9474};
dout[79]={ 16'd13331,-16'd1710,16'd3015,-16'd5065,-16'd8544,16'd9769,16'd9771,16'd3042,-16'd1533,16'd1875,16'd1281,-16'd6350};
dout[80]={ -16'd15224,16'd3247,16'd5006,-16'd1658,16'd6447,-16'd1203,-16'd2511,-16'd8611,-16'd3685,-16'd546,-16'd10492,16'd5665};
dout[81]={ 16'd4318,16'd6926,16'd9647,-16'd3058,16'd4617,16'd1827,16'd5566,-16'd6972,-16'd12811,16'd11271,-16'd9904,16'd5228};
dout[82]={ 16'd2259,16'd3575,16'd5508,-16'd7465,-16'd11076,-16'd2696,-16'd10418,-16'd1549,-16'd7596,-16'd101,16'd10882,-16'd4105};
dout[83]={ -16'd15173,-16'd8289,-16'd4153,-16'd3248,16'd2083,-16'd8824,-16'd4270,-16'd6793,-16'd10723,16'd1123,16'd10853,-16'd6223};
dout[84]={ -16'd5936,16'd6089,16'd7116,16'd9674,-16'd8861,16'd3342,-16'd10828,16'd3441,16'd6225,-16'd815,16'd3252,16'd2240};
dout[85]={ -16'd8147,16'd5039,-16'd9654,-16'd7767,16'd2553,-16'd7980,16'd4736,-16'd5337,16'd751,-16'd9482,16'd11898,16'd4997};
dout[86]={ -16'd1166,-16'd5888,16'd1280,16'd7667,16'd2619,16'd11636,-16'd1945,16'd1375,-16'd4117,16'd8753,-16'd1165,16'd11146};
dout[87]={ 16'd100,16'd9620,16'd8032,-16'd7282,-16'd13759,-16'd4648,-16'd2323,-16'd10309,16'd905,-16'd3167,16'd5564,-16'd3983};
dout[88]={ -16'd17825,-16'd1417,16'd5904,16'd10283,16'd5919,-16'd5557,-16'd11348,-16'd8157,-16'd2027,16'd3896,-16'd6247,16'd12949};
dout[89]={ -16'd9628,16'd5279,16'd11300,16'd1653,16'd2476,16'd823,16'd4932,16'd4759,16'd7045,16'd2599,16'd9766,16'd4500};
dout[90]={ -16'd26059,-16'd2608,16'd6544,16'd13674,16'd7114,16'd5426,16'd3895,-16'd840,-16'd7532,16'd7270,16'd9972,16'd10544};
dout[91]={ -16'd6431,16'd907,16'd12391,16'd5304,-16'd2108,16'd10116,16'd3261,-16'd1717,-16'd225,-16'd6611,16'd3741,-16'd6991};
dout[92]={ 16'd1345,16'd4104,16'd12065,-16'd3992,16'd8188,-16'd7794,16'd6011,-16'd7001,-16'd4439,16'd7094,16'd7798,16'd528};
dout[93]={ 16'd12007,16'd11885,-16'd7319,16'd4404,-16'd9017,16'd477,-16'd8277,-16'd2944,16'd823,16'd6933,16'd7356,16'd4596};
dout[94]={ -16'd5383,-16'd10150,-16'd3602,16'd11115,-16'd5023,-16'd10273,-16'd2175,16'd9559,16'd140,-16'd10763,-16'd117,16'd1714};
dout[95]={ 16'd38887,-16'd3527,16'd4443,16'd2565,-16'd2868,16'd6348,-16'd10153,16'd3552,-16'd13081,-16'd6142,16'd9989,-16'd9608};
dout[96]={ -16'd2706,-16'd4971,16'd2867,16'd376,16'd10536,16'd7485,16'd8181,16'd6500,-16'd7332,-16'd5139,16'd8116,-16'd5390};
dout[97]={ -16'd15343,16'd6204,-16'd1835,-16'd11735,16'd856,16'd5712,16'd11681,16'd10284,-16'd5390,16'd3771,-16'd10452,-16'd10033};
dout[98]={ -16'd2288,16'd11313,16'd6176,-16'd4633,16'd4059,16'd11626,-16'd8901,-16'd13060,16'd7603,16'd7700,16'd5927,-16'd5969};
dout[99]={ 16'd13345,16'd8518,16'd1136,-16'd5964,16'd8640,16'd11951,-16'd4167,-16'd2387,-16'd2890,16'd1541,-16'd7046,-16'd9518};
dout[100]={ 16'd10666,16'd9617,16'd3878,-16'd5802,-16'd8470,16'd9321,-16'd5642,16'd7585,-16'd4252,16'd11439,16'd9263,16'd7784};
dout[101]={ -16'd12484,-16'd6007,-16'd9092,16'd22,16'd387,16'd1912,-16'd9364,16'd865,-16'd4350,-16'd9012,16'd10456,16'd5892};
dout[102]={ -16'd304,-16'd3722,-16'd9202,-16'd4766,16'd8434,-16'd1947,-16'd5139,16'd4949,16'd10327,-16'd9430,-16'd4288,-16'd7285};
dout[103]={ -16'd6946,-16'd1939,-16'd1677,16'd10956,16'd8365,-16'd1867,-16'd10657,-16'd4263,16'd1905,16'd6244,16'd3476,16'd4809};
dout[104]={ 16'd4602,16'd7545,16'd9043,16'd7807,-16'd268,16'd7155,16'd6554,-16'd4544,16'd2396,16'd7335,16'd866,16'd12589};
dout[105]={ -16'd16294,-16'd1390,-16'd8912,-16'd7730,16'd3264,-16'd7584,-16'd2813,-16'd9374,16'd11436,16'd12570,16'd5599,-16'd4140};
dout[106]={ -16'd14640,-16'd6446,16'd6357,16'd903,16'd1718,-16'd8799,16'd5072,-16'd6279,16'd6781,16'd14563,16'd2804,16'd8083};
dout[107]={ 16'd19686,16'd5294,16'd1283,-16'd1490,-16'd14448,-16'd8285,-16'd4491,16'd1201,-16'd1186,16'd4527,-16'd1252,16'd4851};
dout[108]={ 16'd8971,16'd1979,16'd6936,-16'd2413,-16'd11882,-16'd8882,-16'd746,-16'd2529,16'd1034,16'd11507,-16'd7613,16'd3321};
dout[109]={ 16'd6200,16'd10349,16'd12125,16'd2762,-16'd1223,16'd7180,16'd3475,16'd11422,-16'd9987,16'd963,-16'd740,-16'd2319};
dout[110]={ 16'd11483,-16'd10057,-16'd4189,-16'd6134,-16'd97,16'd12801,16'd4031,-16'd9342,-16'd6486,16'd1355,-16'd7764,16'd1534};
dout[111]={ -16'd12423,16'd1389,-16'd12337,16'd575,-16'd3592,16'd253,-16'd2279,16'd12527,-16'd2511,-16'd2002,16'd2113,-16'd72};
dout[112]={ 16'd12385,16'd3253,16'd2745,-16'd1454,16'd2110,16'd5436,-16'd6984,-16'd847,16'd2092,-16'd7084,16'd6859,-16'd3535};
dout[113]={ -16'd16776,-16'd6165,-16'd5641,-16'd280,-16'd3537,-16'd7048,16'd4779,16'd5712,16'd11621,16'd12153,-16'd12112,-16'd8419};
dout[114]={ 16'd25045,-16'd2202,-16'd5828,-16'd13144,16'd7553,16'd4387,-16'd12311,-16'd4076,-16'd5395,16'd8637,16'd5664,-16'd7388};
dout[115]={ -16'd15030,16'd6024,16'd2807,-16'd7604,-16'd6807,16'd3599,16'd10404,16'd10001,16'd2950,-16'd4333,-16'd5619,-16'd5502};
dout[116]={ -16'd5438,-16'd2514,16'd631,-16'd1781,16'd3265,16'd4737,-16'd8315,-16'd9987,-16'd9940,-16'd1586,16'd11541,16'd1201};
dout[117]={ 16'd298,-16'd5046,-16'd6291,-16'd384,16'd10165,16'd9634,16'd10883,-16'd2976,-16'd9393,-16'd6802,-16'd1522,-16'd3150};
dout[118]={ -16'd12337,16'd1475,-16'd7677,-16'd6302,-16'd3450,16'd1033,16'd1138,-16'd1776,16'd5476,-16'd6960,16'd7868,-16'd7076};
dout[119]={ 16'd8087,16'd6636,-16'd5224,-16'd6237,16'd8208,16'd3656,16'd617,16'd9301,16'd6313,16'd757,16'd4633,16'd3899};
dout[120]={ 16'd1548,-16'd7911,16'd9784,16'd7515,16'd2643,16'd7490,16'd8384,-16'd922,16'd6392,-16'd11060,16'd5720,-16'd9063};
dout[121]={ -16'd7919,16'd7579,16'd2092,-16'd3643,-16'd9911,-16'd8284,-16'd10801,-16'd8579,16'd3771,16'd1703,16'd8176,16'd4785};
dout[122]={ -16'd8524,16'd9356,16'd6524,16'd1758,16'd1306,16'd9092,16'd6233,-16'd5628,16'd10911,16'd10214,-16'd1469,16'd81};
dout[123]={ -16'd15784,-16'd1396,-16'd5396,-16'd3316,16'd9989,16'd8519,-16'd4148,-16'd2416,-16'd8896,16'd10421,16'd4109,-16'd3999};
dout[124]={ -16'd16203,16'd8097,16'd2937,-16'd1878,-16'd12458,-16'd6382,16'd8285,16'd1366,-16'd7771,-16'd4238,16'd1690,16'd85};
dout[125]={ 16'd2438,16'd4397,16'd6072,16'd9490,16'd10435,-16'd10454,16'd6666,16'd4891,16'd688,-16'd9668,16'd8998,-16'd8762};
dout[126]={ -16'd6209,16'd10834,16'd10159,-16'd1709,16'd3621,16'd3514,16'd6774,16'd10342,16'd7383,-16'd3110,-16'd4161,-16'd4488};
dout[127]={ -16'd5409,-16'd7689,16'd4929,16'd8754,-16'd8546,-16'd3861,-16'd6005,16'd528,-16'd7169,-16'd9483,-16'd1708,16'd3630};
dout[128]={ -16'd26917,16'd5597,16'd1462,-16'd6495,16'd11881,-16'd5624,-16'd3025,16'd4926,16'd12593,16'd7675,-16'd5973,-16'd3438};
dout[129]={ 16'd4954,-16'd3720,16'd3818,16'd6472,-16'd5992,-16'd8215,16'd10627,-16'd7245,16'd5443,16'd982,16'd2561,16'd12576};
dout[130]={ -16'd24437,-16'd5112,-16'd223,-16'd9329,16'd5165,-16'd1673,16'd8920,-16'd374,-16'd2544,16'd5779,-16'd5487,-16'd6669};
dout[131]={ 16'd6790,-16'd4640,-16'd1283,16'd8491,-16'd6446,-16'd6652,16'd10573,16'd5228,-16'd7829,-16'd6718,-16'd12654,16'd6339};
dout[132]={ -16'd10674,-16'd1058,16'd2648,16'd2296,-16'd7853,16'd7051,16'd1386,-16'd2083,-16'd5654,-16'd5214,16'd4982,16'd7726};
dout[133]={ -16'd9825,-16'd3075,16'd9522,-16'd3933,16'd67,-16'd10441,16'd10373,-16'd9270,16'd3894,16'd5202,-16'd11111,-16'd127};
dout[134]={ -16'd12750,-16'd3763,-16'd9584,-16'd14349,-16'd5245,-16'd10433,-16'd4163,16'd8773,16'd10566,16'd6702,16'd193,-16'd9920};
dout[135]={ -16'd13441,-16'd4774,-16'd301,-16'd166,16'd5550,-16'd4704,-16'd3453,16'd2482,-16'd5560,16'd2972,16'd10520,-16'd9806};
dout[136]={ 16'd12550,-16'd9137,-16'd1386,-16'd1710,16'd8813,-16'd6596,-16'd4909,-16'd4866,-16'd5993,-16'd8878,16'd8928,16'd2998};
dout[137]={ -16'd8014,-16'd10359,16'd11888,-16'd4473,-16'd8094,-16'd6617,16'd9779,-16'd11773,16'd1438,-16'd8778,16'd368,-16'd9498};
dout[138]={ -16'd10679,16'd4095,-16'd1140,16'd16602,-16'd9207,-16'd1300,16'd6250,-16'd6188,16'd1329,-16'd1217,-16'd3482,16'd8408};
dout[139]={ -16'd14671,16'd709,16'd6312,16'd374,16'd9235,-16'd5888,16'd1165,16'd2787,16'd2769,16'd4856,-16'd4677,16'd3724};
dout[140]={ 16'd36294,-16'd5304,16'd8396,16'd2626,-16'd9518,-16'd8455,16'd1851,-16'd8535,16'd10138,-16'd5257,-16'd12439,16'd7127};
dout[141]={ -16'd31908,16'd10822,-16'd5674,16'd10726,16'd495,16'd2632,16'd5350,-16'd6545,16'd8196,-16'd2770,16'd1542,16'd9109};
dout[142]={ -16'd15467,16'd5962,16'd5440,-16'd13760,16'd2120,-16'd3969,16'd494,16'd11405,-16'd1075,-16'd5357,16'd8916,-16'd10463};
dout[143]={ 16'd10443,16'd10699,-16'd5690,-16'd1928,-16'd11529,-16'd426,16'd6545,-16'd7327,-16'd14686,-16'd54,-16'd8884,16'd7552};
end

always @ (posedge clk) begin
  w <= dout[addr];
end


endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */
