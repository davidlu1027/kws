module kernel_0_rom (
    input  wire        [ 10:0] addr,
    input  wire               in_valid,
    input  wire               clk,
    output reg signed [ 575:0] w
  );

reg [575:0] dout [0:1199];


initial begin
dout[0]={ -16'd9311,-16'd1672,16'd1768,16'd4936,-16'd5318,16'd5864,-16'd2636,-16'd1277,16'd7449,-16'd6351,16'd2765,-16'd2330,16'd6109,-16'd865,16'd4934,16'd2058,-16'd217,-16'd5379,16'd1362,-16'd6754,16'd1829,-16'd1676,-16'd4226,-16'd5701,16'd4537,-16'd1599,16'd6636,16'd4009,-16'd6895,16'd4415,16'd2762,-16'd7405,16'd7479,16'd7546,16'd6878,-16'd2917};
dout[1]={ -16'd3598,-16'd863,16'd5240,16'd2794,16'd3539,-16'd397,16'd7527,-16'd986,16'd3427,16'd5123,16'd11717,-16'd3942,16'd1643,-16'd10753,-16'd10984,-16'd5052,-16'd5722,16'd4665,16'd2544,16'd3779,-16'd5289,16'd4066,-16'd343,-16'd1504,-16'd6037,16'd2873,-16'd6627,-16'd5704,16'd5966,-16'd5555,-16'd4265,16'd2911,-16'd1998,16'd4313,16'd5404,-16'd5392};
dout[2]={ 16'd1186,16'd3840,-16'd1270,-16'd428,-16'd2512,-16'd321,16'd4827,16'd6769,-16'd2934,16'd3232,16'd3674,16'd4449,-16'd1193,-16'd2557,-16'd2508,16'd416,16'd3219,-16'd2189,16'd1060,-16'd3905,-16'd2232,16'd5877,-16'd7296,16'd3251,-16'd7981,16'd1243,-16'd6492,-16'd5598,-16'd2872,-16'd1191,16'd2950,-16'd4374,16'd6046,16'd619,-16'd343,-16'd8225};
dout[3]={ -16'd2223,16'd4854,16'd4310,-16'd3601,16'd3612,-16'd3803,-16'd2199,16'd5579,16'd5428,-16'd1483,-16'd6819,16'd1785,-16'd5990,-16'd3132,-16'd7162,-16'd288,-16'd2093,16'd2371,16'd305,-16'd3982,-16'd3009,-16'd5658,-16'd8817,16'd2952,-16'd7799,-16'd4364,-16'd2429,16'd4591,-16'd3097,16'd1838,16'd4472,16'd4350,-16'd7386,-16'd3210,16'd4030,-16'd9208};
dout[4]={ -16'd9095,-16'd2406,16'd8409,-16'd5498,-16'd6487,-16'd2540,16'd3263,-16'd3956,16'd6283,-16'd3665,-16'd5960,-16'd6490,16'd5051,16'd4648,-16'd6080,-16'd4888,16'd1019,16'd4665,16'd1479,-16'd6611,-16'd5380,-16'd3955,16'd2113,-16'd800,16'd48,16'd2886,16'd9678,16'd554,-16'd3673,16'd9350,-16'd4,-16'd3272,-16'd1669,16'd2179,-16'd3560,-16'd2203};
dout[5]={ -16'd4171,-16'd3063,16'd3731,-16'd5285,16'd7224,-16'd6207,16'd1774,16'd3608,-16'd2058,16'd2814,16'd7071,-16'd2588,16'd2653,-16'd4612,-16'd1954,16'd6152,16'd7241,16'd498,-16'd1109,-16'd347,-16'd5599,-16'd3192,-16'd6294,-16'd620,16'd5296,16'd3941,-16'd5968,-16'd3992,-16'd994,-16'd4001,16'd3185,-16'd18,16'd303,-16'd3177,16'd9654,-16'd5290};
dout[6]={ 16'd5534,16'd4080,-16'd2130,16'd4032,-16'd3384,-16'd3949,16'd4148,-16'd1980,16'd4344,-16'd1248,16'd4391,-16'd6606,16'd1060,-16'd7355,16'd2182,16'd1174,16'd3987,-16'd1747,-16'd2064,16'd2096,16'd1261,16'd2563,16'd6566,16'd1879,-16'd6456,16'd340,-16'd2205,-16'd3334,16'd2680,16'd6600,16'd4584,-16'd6227,-16'd3500,16'd5574,16'd5347,16'd443};
dout[7]={ 16'd2684,16'd5833,16'd2954,16'd1823,16'd1944,16'd1543,16'd1625,16'd4278,-16'd7002,16'd5033,-16'd5008,-16'd3081,16'd6873,-16'd1105,16'd8121,-16'd1174,-16'd5424,16'd2142,-16'd2004,-16'd5662,16'd4238,-16'd3989,-16'd5210,-16'd1487,16'd1498,-16'd3862,16'd1105,-16'd1684,-16'd2188,16'd4364,16'd7631,-16'd2977,16'd2431,-16'd4896,16'd30,16'd3079};
dout[8]={ 16'd5869,16'd5788,-16'd657,-16'd2235,16'd785,16'd2026,16'd913,16'd2015,-16'd7728,16'd4717,16'd5066,16'd5974,16'd3055,16'd6251,16'd7526,16'd4419,-16'd3087,16'd4818,16'd8529,-16'd4112,-16'd4565,16'd3312,-16'd6028,16'd5355,-16'd546,16'd3015,-16'd370,16'd6226,-16'd994,-16'd7083,16'd967,-16'd11024,16'd1157,16'd2689,-16'd3438,16'd6837};
dout[9]={ 16'd2701,16'd5123,16'd5009,16'd231,16'd5428,16'd557,16'd1491,16'd4828,-16'd5743,16'd3311,-16'd2920,-16'd2240,-16'd7320,16'd5903,16'd7578,-16'd65,-16'd3546,-16'd5503,-16'd5537,16'd958,16'd3150,-16'd6266,-16'd4783,16'd2703,16'd1188,16'd4483,16'd1741,16'd2492,16'd4356,16'd3715,16'd5628,-16'd10452,-16'd6994,16'd1172,16'd4003,-16'd16};
dout[10]={ -16'd3348,16'd6845,16'd4106,-16'd5856,-16'd4111,-16'd1228,-16'd1395,-16'd6412,16'd4518,-16'd7589,16'd520,16'd4568,16'd1554,-16'd8988,-16'd2447,-16'd1179,-16'd6513,16'd6754,-16'd4064,-16'd8117,-16'd7800,-16'd5627,-16'd6002,-16'd1880,-16'd3205,-16'd334,16'd9639,16'd1577,-16'd4621,16'd4933,-16'd3930,16'd6815,-16'd1148,16'd164,16'd1019,16'd2532};
dout[11]={ 16'd1269,16'd5666,-16'd2103,16'd1179,16'd6519,16'd3786,16'd1200,-16'd7372,-16'd1583,-16'd9616,16'd2238,16'd4104,-16'd4684,16'd1352,-16'd959,16'd3500,16'd158,-16'd6860,-16'd7328,16'd2185,16'd4589,16'd3353,16'd4601,-16'd3083,-16'd2307,-16'd3236,-16'd4270,16'd5665,-16'd1681,16'd318,-16'd6570,16'd12,-16'd320,-16'd2019,-16'd8785,-16'd2418};
dout[12]={ 16'd158,-16'd529,-16'd6787,-16'd5290,-16'd2934,-16'd1619,-16'd5769,16'd522,16'd4059,-16'd4803,16'd5054,16'd316,16'd469,16'd4396,-16'd4253,-16'd6558,-16'd6219,-16'd4689,-16'd1154,-16'd6086,16'd4432,16'd2377,16'd6131,16'd2514,16'd2962,16'd11234,16'd1463,16'd7480,-16'd4514,16'd8069,16'd2743,16'd8876,-16'd8156,16'd9165,16'd1238,16'd2806};
dout[13]={ 16'd997,16'd9174,16'd2528,-16'd3914,16'd1685,16'd1475,16'd3597,16'd6028,16'd4396,-16'd2232,-16'd10630,16'd1774,-16'd8434,-16'd8474,16'd4050,-16'd3184,-16'd3592,-16'd8033,-16'd2712,-16'd8884,16'd5476,-16'd5939,-16'd5228,16'd26,-16'd7072,16'd8239,16'd4027,-16'd1028,-16'd2740,16'd79,16'd6644,-16'd3140,-16'd6470,16'd4412,-16'd746,16'd3541};
dout[14]={ -16'd7688,16'd4354,16'd783,16'd6190,-16'd4035,-16'd6624,16'd307,16'd2492,-16'd8333,16'd1617,-16'd1103,16'd7512,-16'd4961,16'd3840,-16'd2963,16'd386,16'd7964,-16'd4531,-16'd2195,-16'd8051,16'd1633,-16'd1311,-16'd613,-16'd4050,16'd4012,-16'd1381,16'd5660,16'd3357,-16'd5545,16'd3793,-16'd4004,-16'd2194,-16'd652,16'd4670,-16'd783,16'd3405};
dout[15]={ -16'd3271,16'd3347,-16'd466,16'd2940,-16'd748,-16'd785,-16'd1531,16'd5680,-16'd1540,-16'd648,-16'd1536,16'd1708,16'd170,16'd5316,16'd638,-16'd3411,16'd7537,-16'd6802,-16'd7515,16'd5915,-16'd1157,-16'd6043,-16'd687,16'd4948,16'd5242,-16'd5766,16'd2011,-16'd5928,-16'd2887,-16'd1934,16'd2184,16'd1786,-16'd5004,16'd5362,-16'd4805,16'd1321};
dout[16]={ 16'd19,-16'd3954,-16'd2171,-16'd3136,16'd1793,-16'd5463,-16'd3785,-16'd6068,-16'd8301,-16'd5976,16'd1506,-16'd6522,16'd4105,-16'd5098,-16'd385,-16'd2831,16'd2652,-16'd6402,-16'd515,-16'd3354,16'd7251,-16'd5173,-16'd3615,16'd5,-16'd5192,-16'd3683,16'd5563,-16'd60,-16'd1277,16'd4963,16'd2686,16'd2485,-16'd4748,16'd5764,-16'd4397,-16'd4965};
dout[17]={ -16'd618,-16'd4862,16'd3118,-16'd4321,-16'd3506,-16'd1084,-16'd2999,-16'd5254,-16'd4784,-16'd1786,16'd7094,-16'd4306,16'd6592,16'd3573,-16'd1964,16'd3800,-16'd1985,16'd3411,-16'd5270,-16'd6171,-16'd1533,16'd4902,-16'd3405,-16'd2562,16'd2305,-16'd4004,16'd6107,-16'd3120,-16'd4479,16'd460,-16'd2595,-16'd2969,-16'd3948,16'd3691,-16'd4582,16'd3870};
dout[18]={ -16'd5031,16'd7201,16'd4841,16'd6077,16'd5222,16'd6257,16'd5329,-16'd3962,16'd2693,-16'd4108,16'd5563,-16'd7706,16'd2037,-16'd1996,16'd3118,-16'd1285,16'd1229,16'd5823,-16'd2209,16'd7627,-16'd760,-16'd5004,-16'd5707,16'd7995,16'd8059,-16'd5462,16'd24,-16'd3696,16'd6709,16'd7049,-16'd5328,-16'd4575,16'd1859,16'd4595,-16'd4291,16'd7649};
dout[19]={ -16'd5449,16'd5452,16'd6084,16'd10273,16'd3052,-16'd1936,16'd2532,-16'd5472,-16'd5974,16'd7050,-16'd1508,-16'd6064,-16'd2624,16'd3959,-16'd2131,-16'd5862,-16'd468,16'd8007,16'd5913,-16'd3394,16'd8444,-16'd7732,-16'd2608,-16'd5024,16'd5115,16'd4010,-16'd5392,16'd2859,16'd6406,16'd3520,16'd220,-16'd6597,16'd4157,16'd3893,-16'd2325,16'd8097};
dout[20]={ -16'd5879,16'd7234,16'd5192,-16'd6461,16'd278,-16'd6321,-16'd2829,-16'd1648,16'd2341,-16'd1797,16'd6627,-16'd4737,16'd1447,-16'd3912,16'd6222,-16'd2704,16'd65,16'd4964,-16'd6058,-16'd2372,16'd22,16'd6788,-16'd30,16'd5175,-16'd6334,16'd7820,-16'd2107,16'd3662,-16'd11004,16'd1892,16'd7267,16'd4439,-16'd5470,16'd10204,16'd3864,-16'd436};
dout[21]={ 16'd664,-16'd511,-16'd1764,-16'd3800,-16'd3363,-16'd5766,-16'd4588,16'd2061,16'd30,16'd4652,16'd4079,-16'd77,-16'd191,-16'd13238,-16'd5079,-16'd1529,-16'd9634,16'd2272,-16'd2164,16'd3444,16'd6966,-16'd5815,16'd258,-16'd2235,16'd5379,16'd4185,16'd348,16'd4114,-16'd455,16'd3690,-16'd2416,16'd8329,16'd3841,16'd5613,-16'd4727,16'd772};
dout[22]={ -16'd8839,16'd4406,16'd4607,16'd6318,-16'd5531,16'd1155,16'd2739,-16'd7572,16'd3454,-16'd7296,16'd3409,16'd4308,16'd77,-16'd1763,16'd1157,-16'd8253,-16'd3519,16'd2266,-16'd390,16'd3445,-16'd2456,16'd963,16'd5920,16'd2446,-16'd4591,16'd1089,16'd4911,16'd2500,-16'd4951,16'd1851,16'd6213,16'd1910,16'd4439,16'd7070,16'd443,-16'd9202};
dout[23]={ 16'd1159,16'd4920,-16'd1927,16'd2093,-16'd1591,16'd2867,-16'd3033,-16'd7912,16'd3574,16'd7402,-16'd12976,16'd4558,16'd5926,16'd1304,16'd2813,16'd3655,16'd824,16'd2997,-16'd6993,-16'd2508,-16'd3027,-16'd8098,-16'd7364,-16'd5348,-16'd7011,16'd3646,-16'd2243,-16'd508,16'd5574,16'd1579,16'd6082,-16'd6855,-16'd2789,-16'd2688,16'd1500,16'd1552};
dout[24]={ -16'd4368,16'd372,16'd6043,16'd10210,-16'd3981,16'd3816,-16'd9488,16'd6880,-16'd1546,16'd3373,16'd3463,-16'd5503,-16'd5799,-16'd2926,-16'd7644,16'd203,16'd5380,16'd3585,16'd5147,16'd2328,-16'd1638,-16'd1201,-16'd292,16'd2331,16'd5287,-16'd3568,-16'd4536,16'd1987,-16'd9573,-16'd1349,-16'd7047,-16'd5555,16'd7020,-16'd459,16'd6066,16'd5847};
dout[25]={ -16'd6874,-16'd7323,16'd6066,-16'd273,-16'd3487,16'd4777,-16'd302,16'd5416,16'd1534,16'd3903,-16'd420,16'd5321,-16'd1837,-16'd4971,16'd7813,16'd4380,-16'd5545,-16'd2313,16'd347,16'd5341,16'd4196,-16'd4320,16'd4188,-16'd6156,-16'd6269,16'd2222,-16'd1594,-16'd1064,-16'd6661,16'd1343,16'd1139,-16'd7570,-16'd1932,16'd6149,-16'd370,-16'd3921};
dout[26]={ -16'd1300,16'd283,16'd2907,-16'd2929,16'd6400,16'd6918,16'd1652,16'd2742,16'd1216,-16'd6620,16'd2652,16'd5959,16'd3397,16'd3359,-16'd495,-16'd6880,-16'd4204,16'd2630,16'd5063,-16'd146,16'd722,-16'd1782,16'd2368,16'd224,16'd4921,-16'd8131,-16'd6782,-16'd4665,-16'd2197,16'd4036,-16'd5015,-16'd687,-16'd4173,-16'd586,16'd535,16'd6049};
dout[27]={ -16'd4297,-16'd6087,-16'd1116,-16'd5738,16'd1092,-16'd5071,16'd3076,-16'd4588,-16'd4370,16'd6058,16'd7595,16'd2334,-16'd7273,-16'd142,16'd766,-16'd5679,-16'd642,-16'd6037,16'd6785,16'd4792,-16'd3774,-16'd3507,16'd3575,16'd4224,-16'd130,-16'd6547,-16'd5736,-16'd462,-16'd700,16'd605,16'd2796,16'd4535,-16'd6419,16'd5234,-16'd7145,16'd5959};
dout[28]={ 16'd5839,-16'd6124,16'd2562,-16'd4092,16'd7029,-16'd4669,-16'd3830,16'd2127,-16'd3284,16'd8813,-16'd1217,16'd4141,16'd956,16'd2940,-16'd2054,16'd2281,16'd4967,-16'd3823,-16'd4728,-16'd1681,-16'd4398,-16'd6766,16'd1043,-16'd5510,-16'd1358,-16'd6377,-16'd1928,16'd2133,16'd783,-16'd6521,16'd3747,-16'd1173,-16'd6576,16'd5266,16'd5284,-16'd3117};
dout[29]={ 16'd2758,-16'd383,-16'd6478,16'd3360,-16'd3727,-16'd6616,-16'd2098,16'd3006,-16'd1371,-16'd1350,-16'd3296,-16'd7308,16'd6780,16'd2634,16'd1154,16'd3029,16'd4933,16'd677,16'd6812,16'd1419,-16'd2697,16'd4438,-16'd8579,-16'd6657,-16'd7774,-16'd1584,16'd4659,-16'd4142,16'd4328,16'd137,-16'd1785,16'd4891,-16'd6497,-16'd6804,16'd6748,16'd5253};
dout[30]={ -16'd1875,-16'd9166,16'd3069,-16'd2530,16'd340,-16'd5018,-16'd5707,-16'd657,-16'd5745,16'd5858,16'd4869,16'd5390,-16'd727,-16'd13461,16'd8531,-16'd1132,16'd3822,-16'd1365,16'd290,-16'd7886,-16'd893,16'd70,16'd5786,-16'd865,-16'd6196,16'd7892,-16'd2233,16'd4192,-16'd2595,-16'd2147,16'd9719,16'd941,-16'd5974,-16'd361,16'd3220,16'd9197};
dout[31]={ -16'd9241,16'd4883,-16'd1465,-16'd1455,16'd4589,-16'd5345,-16'd9333,-16'd3679,16'd1599,-16'd5880,16'd4413,16'd3171,-16'd6706,-16'd7836,-16'd2987,-16'd489,-16'd5992,-16'd4236,16'd2159,16'd2749,-16'd8193,16'd1657,-16'd4274,-16'd5455,-16'd2846,16'd5329,-16'd1079,-16'd381,16'd657,16'd669,16'd1700,-16'd1274,16'd1531,-16'd3212,16'd3031,-16'd3193};
dout[32]={ -16'd7243,-16'd6507,16'd4066,-16'd6228,-16'd1567,-16'd7439,-16'd4897,-16'd3211,-16'd8702,-16'd7899,-16'd1871,16'd7482,-16'd4503,-16'd4240,16'd469,-16'd4489,-16'd6958,16'd1601,-16'd2804,-16'd7687,-16'd4107,16'd1536,16'd439,16'd3873,16'd6315,-16'd3377,-16'd5676,-16'd88,-16'd3087,16'd708,16'd1681,-16'd898,-16'd4457,16'd648,-16'd7742,-16'd3695};
dout[33]={ 16'd4142,16'd4298,16'd3788,16'd3022,-16'd73,16'd924,-16'd8099,16'd3456,-16'd4965,-16'd2139,-16'd6823,16'd5402,16'd1253,16'd909,-16'd3858,16'd4404,16'd4247,16'd2721,16'd2809,-16'd4693,-16'd4707,16'd2859,16'd3472,-16'd5806,-16'd1962,16'd5775,16'd3830,16'd549,16'd2808,16'd7678,16'd2064,-16'd5228,-16'd6544,-16'd4577,-16'd2596,-16'd2631};
dout[34]={ 16'd758,-16'd4027,16'd6587,-16'd3715,-16'd6614,-16'd969,16'd2202,-16'd1903,-16'd4676,-16'd2401,-16'd3177,-16'd1409,16'd7469,16'd4614,16'd391,16'd1345,16'd154,-16'd150,-16'd127,16'd746,-16'd2130,-16'd1039,-16'd2687,16'd451,-16'd6723,-16'd1147,-16'd3931,-16'd4514,-16'd9236,-16'd3755,16'd3951,16'd6290,-16'd7179,16'd1906,-16'd897,16'd3373};
dout[35]={ -16'd88,16'd3597,16'd3414,-16'd2838,-16'd7691,16'd2874,16'd4664,-16'd6820,16'd4196,16'd3205,-16'd5063,-16'd2039,-16'd1960,-16'd3089,-16'd1896,-16'd1303,16'd7133,-16'd4067,16'd4396,16'd899,16'd1124,16'd3403,16'd5028,16'd5640,16'd5470,-16'd772,-16'd3913,16'd4579,-16'd4301,16'd6526,16'd3656,-16'd4745,-16'd3519,16'd2825,16'd472,-16'd152};
dout[36]={ 16'd4440,16'd2632,16'd3360,-16'd1232,16'd4583,-16'd4745,16'd2979,16'd5349,16'd3328,16'd1076,16'd213,-16'd2963,-16'd5700,16'd3590,-16'd3264,-16'd5094,-16'd5435,-16'd5491,-16'd3332,-16'd6732,16'd1707,16'd3327,16'd5298,-16'd6596,-16'd7751,16'd6773,16'd481,16'd1592,-16'd6165,16'd406,-16'd477,16'd6984,-16'd8141,16'd8405,16'd6251,-16'd4094};
dout[37]={ 16'd36,-16'd1907,16'd2584,16'd2222,16'd4436,-16'd3900,16'd6837,-16'd5100,16'd1747,-16'd4853,16'd4240,-16'd111,-16'd3165,-16'd2648,-16'd3209,-16'd76,16'd363,-16'd233,-16'd3300,-16'd5494,-16'd1953,16'd4789,16'd3741,16'd3204,-16'd2940,-16'd1290,-16'd549,16'd3090,16'd2191,-16'd2436,-16'd9020,16'd1489,-16'd7329,-16'd4079,16'd3578,16'd3374};
dout[38]={ -16'd5653,-16'd7149,-16'd2805,16'd6087,16'd3548,16'd4983,-16'd6033,-16'd441,16'd2415,-16'd4037,16'd6385,-16'd695,-16'd5884,-16'd2499,-16'd4304,16'd926,-16'd5129,16'd3518,16'd8069,-16'd3554,16'd6717,16'd2057,16'd3610,-16'd2803,-16'd2623,-16'd6633,16'd2874,16'd3135,16'd5537,-16'd6113,16'd555,-16'd2355,16'd2976,16'd5263,-16'd5998,16'd8661};
dout[39]={ 16'd2507,-16'd1030,16'd3025,16'd4819,-16'd4193,-16'd5282,-16'd3926,-16'd2475,16'd2285,16'd553,16'd1084,-16'd8125,16'd3895,16'd1271,-16'd3742,-16'd4184,-16'd5294,16'd4142,-16'd5400,-16'd3809,-16'd5516,16'd5486,-16'd1495,-16'd1135,16'd1604,16'd3854,16'd6135,16'd1349,16'd7056,16'd636,-16'd1596,-16'd2875,-16'd1241,16'd3495,16'd865,16'd8850};
dout[40]={ 16'd1026,-16'd5755,16'd4161,-16'd9383,-16'd8651,16'd1970,16'd3153,-16'd4652,-16'd5945,-16'd2509,-16'd8629,-16'd3724,16'd4139,-16'd13765,16'd2981,16'd1555,16'd3473,-16'd646,16'd4468,-16'd7470,16'd1610,16'd544,16'd1158,-16'd3104,-16'd446,-16'd2834,-16'd10386,-16'd1881,16'd2087,-16'd4399,16'd469,16'd5288,-16'd4615,16'd1716,-16'd6970,16'd4084};
dout[41]={ -16'd9584,-16'd4142,-16'd8080,16'd255,-16'd2528,16'd6314,-16'd10030,-16'd4434,-16'd3753,-16'd4349,-16'd828,-16'd1960,16'd1258,-16'd4743,16'd1621,-16'd8444,-16'd1911,16'd2374,-16'd3471,-16'd5694,-16'd5586,16'd6856,16'd6954,-16'd7200,16'd4504,-16'd1824,-16'd4507,-16'd3912,-16'd275,16'd1153,-16'd120,-16'd1805,-16'd8048,-16'd2758,-16'd5613,-16'd1890};
dout[42]={ -16'd3221,-16'd226,16'd7339,16'd3650,16'd726,16'd1241,-16'd8552,16'd1597,16'd2987,16'd3682,-16'd442,-16'd2205,-16'd412,-16'd8435,16'd8473,-16'd1660,-16'd7534,16'd1627,16'd598,-16'd3471,-16'd2636,16'd273,-16'd1823,-16'd2790,16'd2412,-16'd3664,-16'd6693,-16'd3542,16'd4963,-16'd8919,16'd6791,16'd2830,-16'd9461,16'd270,16'd215,-16'd5428};
dout[43]={ -16'd5654,-16'd2769,-16'd1003,16'd5022,16'd3823,-16'd7855,16'd2140,-16'd7153,-16'd2393,16'd4545,-16'd10961,-16'd5983,-16'd3207,-16'd2773,16'd7038,-16'd8322,16'd959,-16'd2525,-16'd6396,16'd2635,16'd4589,-16'd6110,16'd3617,-16'd2093,16'd4298,16'd8715,-16'd6926,-16'd6556,-16'd6407,-16'd1464,-16'd5278,-16'd5358,16'd1609,16'd8034,-16'd4774,16'd10039};
dout[44]={ -16'd4960,16'd2928,16'd943,16'd3577,-16'd7176,-16'd6026,-16'd4579,-16'd2471,-16'd5739,16'd558,-16'd103,16'd150,16'd2157,-16'd2806,16'd6746,-16'd1218,-16'd2102,-16'd5559,-16'd5553,-16'd6304,-16'd1810,-16'd2907,-16'd1469,16'd6809,-16'd1703,16'd5986,-16'd1582,16'd332,16'd5256,16'd2496,-16'd4999,-16'd2494,16'd3366,-16'd6144,-16'd2163,-16'd1722};
dout[45]={ -16'd4949,-16'd3067,-16'd1363,-16'd1454,-16'd1848,-16'd1503,-16'd1701,16'd3258,16'd2768,16'd3816,-16'd433,16'd6203,16'd2349,16'd3591,16'd2181,-16'd2761,16'd1921,-16'd3745,-16'd4837,16'd2922,-16'd6247,16'd8450,-16'd413,16'd563,16'd3651,16'd5907,16'd6440,-16'd8529,16'd276,16'd4514,16'd2958,16'd4824,-16'd2501,16'd2608,-16'd6144,16'd4053};
dout[46]={ 16'd1307,16'd139,-16'd36,-16'd5210,-16'd869,-16'd6186,-16'd4635,16'd3410,-16'd708,-16'd910,16'd2540,-16'd3254,16'd2234,16'd6438,16'd3846,-16'd8162,-16'd5457,16'd3702,-16'd4191,16'd3563,16'd4720,16'd1407,16'd5330,16'd2326,16'd212,-16'd6146,-16'd1986,-16'd599,-16'd4553,-16'd2,16'd2072,-16'd5316,-16'd5377,16'd1271,-16'd2915,16'd2703};
dout[47]={ 16'd4030,16'd630,-16'd5980,-16'd2216,16'd1746,-16'd219,-16'd5197,16'd2588,-16'd6746,-16'd4437,-16'd7642,16'd4422,-16'd905,16'd4425,-16'd358,-16'd8255,16'd3262,-16'd4977,-16'd1659,16'd2717,16'd7946,16'd1271,16'd3954,-16'd2533,-16'd2952,-16'd7004,-16'd1280,-16'd5761,16'd7204,-16'd3366,16'd3107,-16'd3781,16'd6207,16'd9099,-16'd5841,16'd4382};
dout[48]={ 16'd7030,-16'd5528,-16'd2469,16'd4989,16'd742,16'd894,16'd6822,-16'd1736,16'd6185,16'd5931,-16'd4256,16'd3538,16'd4671,16'd5149,-16'd4964,16'd3502,16'd6159,16'd5181,-16'd465,16'd3233,16'd168,16'd5200,16'd1778,-16'd569,16'd3011,16'd3360,16'd6359,16'd4599,16'd302,-16'd2147,-16'd7777,-16'd4880,16'd1714,16'd550,16'd3001,16'd1904};
dout[49]={ -16'd5776,-16'd794,-16'd2290,16'd7239,-16'd4379,16'd543,-16'd4388,16'd5602,16'd2693,16'd4859,16'd6177,-16'd5168,16'd4722,16'd1869,16'd6233,16'd2707,16'd4999,16'd1442,16'd8082,-16'd5958,-16'd114,-16'd7867,16'd5078,-16'd2097,-16'd10598,16'd3778,16'd7537,16'd1037,-16'd4030,16'd4483,16'd731,-16'd729,16'd2320,-16'd5827,16'd137,16'd3338};
dout[50]={ -16'd5662,16'd1445,-16'd2633,16'd5555,16'd3842,-16'd4864,16'd1585,16'd1587,-16'd5874,-16'd3526,-16'd5816,16'd1101,16'd6454,-16'd8049,16'd5362,-16'd3607,16'd2701,16'd1391,16'd3561,-16'd8343,16'd2627,16'd7662,-16'd2150,16'd4073,16'd2060,-16'd4841,-16'd10267,-16'd6406,-16'd499,16'd820,16'd6091,16'd5317,16'd2154,16'd1489,16'd7397,16'd7372};
dout[51]={ -16'd3272,-16'd4740,-16'd3091,-16'd6517,-16'd2552,16'd2092,-16'd6404,16'd2979,16'd5672,16'd2320,16'd5185,-16'd1449,16'd6739,-16'd3682,16'd1422,-16'd3621,-16'd544,16'd1027,16'd3070,16'd4268,16'd3138,-16'd7111,16'd6083,-16'd10890,16'd341,16'd1823,-16'd6847,16'd4477,-16'd5301,-16'd5718,16'd5980,-16'd5304,16'd4435,16'd3565,16'd1036,16'd1232};
dout[52]={ 16'd1679,16'd2420,-16'd3602,16'd6538,16'd2413,-16'd480,16'd3331,-16'd6179,-16'd8502,-16'd6264,16'd7092,-16'd4337,-16'd5633,-16'd10738,-16'd5682,16'd1809,-16'd1964,16'd2715,16'd2457,16'd2776,16'd865,-16'd1232,16'd333,16'd3238,-16'd2138,-16'd5564,-16'd11472,16'd5558,-16'd499,-16'd8440,16'd4159,16'd3276,16'd282,-16'd2717,16'd2594,16'd73};
dout[53]={ -16'd5970,16'd7610,16'd8788,16'd5085,-16'd3517,-16'd7602,-16'd5552,-16'd2092,16'd4795,-16'd2128,-16'd5271,-16'd2437,16'd4615,-16'd699,16'd7848,-16'd4857,16'd7997,16'd3155,16'd4940,-16'd6744,-16'd2962,-16'd94,-16'd3604,-16'd4492,16'd1077,16'd5874,16'd1787,-16'd6993,-16'd7379,-16'd1002,-16'd6701,16'd2361,-16'd7144,-16'd667,-16'd621,-16'd1495};
dout[54]={ -16'd5934,16'd5096,-16'd2824,-16'd3151,-16'd4298,16'd5202,-16'd5910,-16'd8982,-16'd3285,-16'd4252,16'd3555,-16'd6166,16'd6813,16'd1246,16'd6030,16'd3635,16'd8297,16'd4284,16'd3046,-16'd6370,-16'd963,16'd2879,-16'd3003,-16'd633,16'd5706,16'd5869,-16'd7136,-16'd4296,-16'd2190,-16'd2854,16'd2678,-16'd6193,-16'd8409,16'd3052,16'd1564,16'd3737};
dout[55]={ -16'd3446,16'd3187,16'd3724,16'd6988,16'd1550,16'd5335,16'd5764,-16'd5664,-16'd3037,16'd6145,16'd6539,16'd5574,16'd2521,16'd4657,16'd1863,16'd3775,-16'd807,-16'd629,16'd1161,16'd1938,-16'd377,16'd3396,-16'd2618,16'd1996,-16'd5753,16'd2530,-16'd2779,16'd4811,16'd46,-16'd5580,-16'd4084,-16'd314,-16'd4979,16'd3694,-16'd1832,-16'd2715};
dout[56]={ 16'd3065,-16'd6875,-16'd5032,16'd3416,16'd5489,16'd1279,-16'd5695,-16'd6169,16'd3081,16'd2274,-16'd804,16'd3546,-16'd261,16'd6354,16'd3101,16'd4958,16'd1099,-16'd4747,-16'd3979,16'd5504,-16'd6603,-16'd7282,-16'd5802,-16'd2445,-16'd6439,-16'd3075,-16'd2751,-16'd7903,16'd702,16'd3031,-16'd4353,16'd3692,16'd874,16'd4977,16'd4655,-16'd2752};
dout[57]={ 16'd2620,-16'd6733,16'd1289,16'd6125,-16'd3810,-16'd1162,-16'd6293,16'd6882,-16'd3067,16'd4997,16'd1404,16'd4377,16'd1292,-16'd6777,-16'd379,16'd1907,16'd7546,-16'd566,-16'd3295,-16'd4471,-16'd4309,16'd5752,16'd3742,-16'd4427,-16'd8510,-16'd622,16'd6889,16'd455,-16'd2742,-16'd5027,-16'd754,-16'd8905,-16'd354,16'd7122,16'd3962,16'd6287};
dout[58]={ 16'd803,16'd4721,16'd5627,16'd4885,-16'd4340,16'd6327,-16'd5702,16'd3509,-16'd4166,-16'd541,-16'd3018,-16'd6364,-16'd5966,-16'd2706,16'd835,-16'd3759,-16'd4307,16'd439,-16'd5474,16'd1879,-16'd4514,-16'd7143,-16'd6815,16'd5204,-16'd2194,16'd2200,16'd4837,-16'd7779,16'd6999,16'd1585,16'd5687,-16'd7427,-16'd696,-16'd3365,-16'd8565,16'd6381};
dout[59]={ 16'd473,-16'd4262,16'd59,-16'd3603,16'd6488,16'd4917,-16'd3319,-16'd2772,-16'd5147,-16'd399,-16'd3344,16'd5818,-16'd7183,-16'd908,-16'd4357,-16'd2530,16'd715,-16'd765,-16'd234,16'd7549,-16'd4385,16'd1128,16'd1643,-16'd6089,16'd775,-16'd5762,16'd8917,16'd2796,16'd4506,-16'd2584,-16'd1389,16'd6021,16'd5140,16'd47,16'd6263,16'd3617};
dout[60]={ -16'd4364,16'd2562,-16'd3070,-16'd4771,-16'd2331,16'd2350,16'd6693,16'd4110,16'd4733,-16'd6210,-16'd231,-16'd3002,16'd6126,16'd137,16'd7103,-16'd5927,-16'd5079,16'd1701,-16'd5429,-16'd4765,-16'd4234,16'd6709,-16'd6138,-16'd205,-16'd2648,-16'd5702,16'd6077,-16'd4356,16'd927,-16'd7162,16'd5663,16'd9996,-16'd4356,-16'd3784,16'd4227,16'd8396};
dout[61]={ -16'd4661,16'd6282,16'd3599,-16'd337,16'd1063,16'd7404,16'd6704,-16'd4425,16'd2058,-16'd1030,16'd619,16'd1714,-16'd2251,-16'd5839,16'd8479,-16'd147,-16'd7496,-16'd6245,-16'd385,16'd1210,-16'd2951,-16'd3380,16'd122,-16'd6307,16'd328,16'd7658,16'd108,-16'd3998,-16'd7078,-16'd7008,16'd3818,-16'd1315,-16'd661,16'd1197,-16'd6675,16'd16};
dout[62]={ -16'd11582,16'd1567,16'd3176,-16'd2976,-16'd1758,16'd1817,-16'd1983,16'd2568,-16'd909,-16'd4867,16'd7060,-16'd7029,-16'd2198,-16'd10707,-16'd349,-16'd8942,-16'd9309,-16'd4274,-16'd1723,16'd5550,16'd1368,-16'd8390,16'd2728,16'd2606,16'd1333,-16'd4379,-16'd9356,-16'd1519,16'd929,-16'd6092,-16'd1610,16'd4657,-16'd1469,16'd836,16'd7045,-16'd3489};
dout[63]={ -16'd2526,-16'd4508,16'd7422,16'd5695,-16'd5502,16'd5211,16'd141,-16'd4585,16'd2961,-16'd497,16'd3077,-16'd2656,-16'd2492,-16'd6450,16'd4644,16'd1299,16'd3124,-16'd1287,-16'd3588,16'd5234,-16'd3066,-16'd2479,16'd3741,-16'd759,-16'd2427,-16'd3570,-16'd4600,16'd7179,-16'd3000,16'd4646,-16'd9083,16'd3617,-16'd4079,16'd1227,-16'd1678,16'd7198};
dout[64]={ -16'd9256,-16'd841,16'd3168,16'd342,-16'd5665,16'd5929,-16'd1634,-16'd2764,-16'd5587,-16'd5968,-16'd2924,16'd7383,-16'd4679,16'd3029,16'd6313,16'd1185,-16'd5536,16'd5092,16'd2990,-16'd7390,-16'd5134,16'd4366,16'd2441,-16'd6153,-16'd5000,16'd6672,-16'd4574,16'd1830,16'd5633,16'd284,-16'd8753,-16'd1721,-16'd2975,16'd2999,-16'd1770,16'd3046};
dout[65]={ -16'd3424,-16'd8404,-16'd6445,16'd688,-16'd7268,16'd1504,16'd3472,-16'd1234,16'd1154,16'd4187,-16'd4343,-16'd3172,16'd991,16'd297,-16'd2255,16'd4005,-16'd3579,16'd7176,16'd3286,-16'd3271,-16'd3566,16'd5763,16'd620,-16'd2920,-16'd3524,16'd6008,-16'd4812,-16'd5370,-16'd1505,-16'd3448,16'd2594,16'd6113,-16'd1840,16'd7528,-16'd6490,16'd6394};
dout[66]={ 16'd2297,-16'd2924,-16'd356,-16'd7374,16'd5483,16'd2365,-16'd3615,-16'd7385,16'd2096,-16'd2329,-16'd1670,16'd8091,16'd4687,-16'd5031,-16'd3929,16'd1032,-16'd5183,16'd1702,-16'd3570,16'd1262,-16'd6036,16'd1922,-16'd1360,16'd5861,-16'd7834,16'd5807,-16'd4978,-16'd2271,16'd5149,16'd6555,-16'd3934,16'd3119,16'd3439,-16'd2716,16'd5367,16'd100};
dout[67]={ -16'd6364,-16'd6857,-16'd6674,16'd3916,-16'd100,-16'd2801,16'd8053,-16'd6065,16'd5173,16'd684,-16'd4090,16'd6072,-16'd4565,-16'd2142,16'd4342,-16'd1957,16'd4079,-16'd289,16'd7451,-16'd7191,16'd1505,16'd888,-16'd3583,-16'd4685,16'd270,16'd4757,-16'd2234,16'd4749,16'd2802,-16'd1095,-16'd3846,16'd533,-16'd5726,16'd1141,-16'd7352,16'd1400};
dout[68]={ 16'd6720,16'd778,-16'd4245,-16'd2357,-16'd1830,16'd4364,-16'd757,-16'd6311,-16'd7003,16'd5802,16'd5094,-16'd6210,-16'd4251,-16'd2691,16'd5920,16'd2746,-16'd2561,16'd4230,-16'd1426,-16'd3328,16'd9704,-16'd512,-16'd5916,-16'd5705,-16'd11039,-16'd4582,16'd3875,-16'd219,16'd3160,-16'd3863,-16'd5182,16'd667,-16'd67,16'd8875,-16'd186,-16'd469};
dout[69]={ -16'd1634,-16'd3336,16'd871,-16'd3159,-16'd8154,-16'd1524,-16'd5382,16'd2432,-16'd6312,-16'd1057,16'd7046,-16'd5486,16'd628,16'd1936,-16'd6861,16'd6355,-16'd5200,-16'd1591,16'd2650,16'd851,16'd3388,-16'd9262,-16'd5384,-16'd6736,-16'd943,16'd128,16'd1361,16'd4182,-16'd5404,-16'd2807,-16'd3655,16'd2353,-16'd5513,-16'd2085,-16'd4458,16'd3967};
dout[70]={ 16'd10828,16'd4413,-16'd925,-16'd3017,16'd2750,16'd4481,-16'd4747,-16'd604,16'd2425,-16'd5094,16'd2799,-16'd9621,-16'd8940,-16'd2212,-16'd9113,-16'd2853,16'd2358,-16'd3567,-16'd9690,16'd1176,-16'd6170,-16'd845,-16'd13415,-16'd4159,-16'd1300,16'd2236,-16'd573,16'd6685,-16'd1150,-16'd1120,16'd8231,16'd6506,-16'd1797,16'd2443,-16'd867,16'd5216};
dout[71]={ 16'd5105,16'd2610,16'd5281,-16'd4281,16'd80,16'd707,16'd1423,-16'd2147,-16'd8389,-16'd7752,16'd6509,-16'd1843,16'd3081,-16'd3321,16'd6928,16'd5467,-16'd9361,-16'd7205,-16'd8756,16'd3060,16'd4824,16'd5269,16'd2196,-16'd6511,-16'd4669,-16'd1975,-16'd1260,16'd1859,16'd2958,16'd78,16'd8757,16'd6133,-16'd3945,16'd2018,16'd4497,16'd5528};
dout[72]={ 16'd4301,16'd9863,16'd8262,16'd3232,-16'd771,16'd1618,16'd7238,16'd8762,16'd1988,16'd3279,16'd10649,16'd2696,-16'd5237,-16'd1519,-16'd741,-16'd8131,16'd2483,16'd1046,-16'd2076,16'd5705,16'd4944,-16'd1967,16'd7523,-16'd60,-16'd1109,-16'd7447,-16'd6169,-16'd6023,-16'd6113,-16'd6397,-16'd4084,16'd2429,16'd1867,-16'd7990,-16'd6420,16'd1836};
dout[73]={ 16'd1714,-16'd206,-16'd7991,16'd410,-16'd106,-16'd3252,-16'd4937,16'd2836,-16'd3447,-16'd7167,16'd424,16'd2733,-16'd5323,-16'd2344,16'd8314,16'd5485,-16'd2783,-16'd720,16'd1091,16'd764,-16'd1078,16'd5802,-16'd3917,16'd1815,16'd5309,16'd736,16'd5749,-16'd2185,-16'd4378,-16'd1998,-16'd330,-16'd268,-16'd264,16'd6604,-16'd5909,16'd4269};
dout[74]={ 16'd1612,16'd4336,16'd3076,16'd6039,-16'd6672,-16'd1839,-16'd5748,-16'd5108,-16'd2403,16'd2873,-16'd4071,16'd5774,16'd2487,16'd1029,-16'd1313,16'd5282,16'd2330,-16'd646,-16'd2035,16'd5158,16'd2963,-16'd2053,16'd2372,-16'd5348,-16'd1131,-16'd1590,-16'd1975,-16'd1259,-16'd5295,16'd2989,-16'd6725,-16'd886,16'd832,-16'd1351,16'd1616,-16'd759};
dout[75]={ -16'd383,-16'd96,16'd3519,16'd7103,-16'd7183,-16'd449,16'd211,-16'd9169,-16'd365,-16'd979,16'd7323,-16'd4220,-16'd6606,16'd5434,16'd2313,-16'd1682,-16'd1697,16'd696,-16'd9775,16'd217,-16'd1586,16'd4855,16'd4781,-16'd7462,16'd5785,16'd3748,-16'd125,-16'd2716,-16'd3457,16'd6095,16'd3808,-16'd2649,-16'd6645,16'd2491,16'd1474,16'd6732};
dout[76]={ 16'd6250,-16'd6250,-16'd4143,16'd6268,16'd3505,16'd3654,-16'd5590,-16'd2455,-16'd1234,16'd3024,16'd6145,16'd4339,-16'd7394,16'd2543,16'd24,16'd1900,16'd3554,16'd219,16'd196,-16'd1305,16'd538,16'd2280,-16'd7687,-16'd1207,16'd3415,-16'd2422,16'd2775,16'd3158,-16'd3649,16'd1928,16'd1092,-16'd2285,16'd5897,16'd6259,16'd1707,-16'd2962};
dout[77]={ 16'd5456,-16'd5711,-16'd6598,16'd1505,-16'd3450,-16'd6853,16'd2639,-16'd4915,16'd3727,-16'd6761,16'd4321,-16'd2810,16'd3455,-16'd2358,-16'd2982,-16'd4489,16'd11,-16'd9124,-16'd2142,-16'd265,16'd750,-16'd2713,-16'd8172,16'd5098,16'd772,-16'd3369,16'd881,-16'd4881,16'd6264,-16'd4281,-16'd3896,-16'd380,-16'd2452,16'd2047,-16'd5797,16'd5331};
dout[78]={ -16'd992,-16'd5165,-16'd7372,-16'd3340,-16'd7676,16'd4713,16'd3187,16'd4315,-16'd4882,-16'd4833,16'd4935,-16'd2595,16'd5291,16'd6074,16'd4584,-16'd3110,-16'd565,-16'd674,-16'd2909,-16'd3369,16'd1845,16'd410,16'd3948,16'd1840,-16'd6462,16'd3391,16'd2009,16'd5409,-16'd2528,16'd1333,-16'd3323,-16'd2610,-16'd6047,16'd1039,-16'd2529,-16'd508};
dout[79]={ -16'd2146,16'd1579,16'd3045,16'd257,16'd90,-16'd2559,-16'd1553,16'd5958,16'd1220,16'd1819,-16'd1207,-16'd829,16'd3665,16'd4766,-16'd1440,16'd6928,-16'd1531,16'd1865,-16'd2582,16'd6312,16'd5004,16'd2089,16'd5406,16'd8032,-16'd226,16'd2472,16'd1961,-16'd4795,-16'd3617,16'd2354,16'd3203,16'd2824,16'd2862,-16'd279,-16'd6577,-16'd7352};
dout[80]={ 16'd7015,-16'd3515,-16'd21,16'd5963,-16'd878,16'd1605,16'd3650,16'd3336,16'd5541,16'd2799,-16'd2187,-16'd1701,-16'd8812,-16'd8082,-16'd4650,-16'd114,-16'd12381,-16'd625,16'd679,-16'd5091,-16'd5157,-16'd6320,-16'd5819,16'd1687,-16'd478,-16'd857,16'd4133,-16'd919,-16'd681,-16'd849,-16'd1793,16'd459,-16'd10018,-16'd4484,-16'd8602,16'd6912};
dout[81]={ 16'd2092,16'd6983,16'd3934,16'd2775,-16'd2730,-16'd3173,16'd7040,16'd3596,-16'd4569,-16'd9864,16'd4158,-16'd10877,-16'd1949,-16'd13059,16'd4246,16'd1818,-16'd3460,16'd1220,16'd3061,16'd2991,-16'd8922,16'd3215,16'd6241,-16'd5043,-16'd4753,-16'd9328,16'd1688,-16'd2945,-16'd7228,-16'd1156,16'd650,16'd149,-16'd7055,-16'd197,-16'd940,-16'd3977};
dout[82]={ 16'd346,-16'd6381,16'd5782,16'd4463,-16'd7399,-16'd238,-16'd200,16'd7967,16'd3088,-16'd6612,-16'd153,16'd3168,-16'd6222,-16'd6701,-16'd5593,-16'd2290,-16'd7912,-16'd39,-16'd5592,-16'd4618,-16'd6564,16'd7273,16'd3382,-16'd6608,-16'd2159,-16'd11758,-16'd144,-16'd592,-16'd5403,16'd9321,-16'd4614,16'd4376,-16'd7820,-16'd7782,-16'd2571,16'd9423};
dout[83]={ 16'd3665,-16'd1627,-16'd1557,16'd4700,-16'd3902,16'd50,-16'd5861,-16'd4536,16'd1427,16'd1839,16'd4355,-16'd7904,16'd796,-16'd1592,16'd2893,16'd5904,16'd2795,16'd1284,-16'd4278,-16'd4902,-16'd1004,-16'd536,-16'd4026,-16'd1975,16'd2320,16'd3170,-16'd4719,16'd684,-16'd1540,16'd1583,-16'd9524,-16'd6625,16'd1259,-16'd1393,-16'd3248,16'd10056};
dout[84]={ -16'd7163,16'd4483,-16'd4965,-16'd7387,-16'd4781,16'd1291,16'd5370,16'd16,-16'd4989,-16'd3014,-16'd3652,16'd2199,-16'd6088,16'd209,-16'd7408,16'd5087,16'd2471,16'd345,-16'd2703,16'd9067,-16'd7293,-16'd3450,-16'd786,-16'd795,-16'd5201,16'd8546,16'd415,-16'd3639,-16'd2562,-16'd2480,-16'd10974,16'd1017,-16'd3985,16'd1200,16'd3562,16'd4063};
dout[85]={ 16'd6506,16'd4086,-16'd6123,-16'd1758,16'd2931,16'd5161,16'd3810,16'd2189,-16'd1313,-16'd917,-16'd3845,16'd4975,-16'd3272,-16'd7935,-16'd1028,16'd2559,16'd906,16'd4460,-16'd916,-16'd2877,-16'd5707,16'd4070,-16'd2892,-16'd377,-16'd3766,-16'd1313,16'd1433,16'd3855,-16'd6565,-16'd2956,-16'd934,16'd2399,-16'd4382,16'd281,16'd1946,-16'd3307};
dout[86]={ -16'd3537,16'd5922,16'd2494,16'd2195,-16'd101,16'd1562,-16'd3660,-16'd5631,-16'd8319,16'd4359,16'd4178,-16'd4278,16'd4206,16'd4467,-16'd2493,-16'd762,-16'd1141,-16'd8972,-16'd3294,-16'd5685,16'd2623,-16'd1056,-16'd2247,-16'd3461,-16'd6983,16'd5926,16'd5753,16'd2072,-16'd1328,-16'd2025,-16'd5595,-16'd954,-16'd4869,16'd7446,16'd73,-16'd713};
dout[87]={ -16'd3716,16'd2273,-16'd1922,-16'd1352,-16'd5808,-16'd3157,-16'd1877,16'd402,-16'd2578,16'd1715,-16'd7030,16'd5252,16'd3752,16'd1035,16'd27,-16'd3295,16'd3978,16'd4334,-16'd4839,-16'd1762,16'd7104,-16'd6963,16'd5745,16'd3444,16'd4903,-16'd1633,-16'd3315,-16'd3874,-16'd5415,-16'd2031,-16'd3059,16'd5108,-16'd1551,-16'd3324,-16'd8771,-16'd5093};
dout[88]={ 16'd6294,-16'd158,16'd5638,16'd1124,16'd3641,-16'd2916,16'd4875,-16'd2298,-16'd4893,-16'd3854,16'd2174,-16'd2983,-16'd5674,-16'd8010,16'd257,16'd798,16'd6150,-16'd1635,-16'd3458,16'd3666,16'd4658,-16'd3422,-16'd3582,16'd2154,-16'd1455,-16'd3387,16'd1252,16'd4618,16'd3096,16'd4598,-16'd6613,-16'd6685,16'd4522,16'd1068,16'd5614,16'd699};
dout[89]={ -16'd2053,16'd2724,16'd2929,-16'd5437,-16'd385,-16'd868,16'd4807,-16'd4091,16'd1065,-16'd871,16'd2961,-16'd6804,16'd3729,-16'd2455,16'd3002,-16'd670,-16'd6117,-16'd1036,-16'd7440,-16'd1503,-16'd1421,-16'd6663,16'd6309,-16'd134,16'd4043,16'd6221,16'd1175,16'd676,16'd8868,16'd6478,16'd3192,-16'd3753,16'd2427,-16'd5523,-16'd5567,16'd663};
dout[90]={ 16'd924,16'd6291,-16'd5209,16'd1059,-16'd6562,-16'd2390,-16'd2872,16'd4360,-16'd6574,-16'd1276,-16'd5882,16'd2616,-16'd1557,-16'd4974,-16'd6632,-16'd411,-16'd7097,-16'd78,-16'd2029,-16'd5955,-16'd4146,16'd1167,-16'd2284,16'd2523,16'd2550,16'd7875,16'd8132,16'd5909,-16'd5169,-16'd204,-16'd5249,-16'd5074,-16'd218,-16'd509,-16'd4414,16'd5992};
dout[91]={ -16'd5537,-16'd3532,-16'd7001,16'd5615,-16'd3029,-16'd3638,-16'd7484,-16'd1291,-16'd6008,16'd2185,-16'd7898,16'd3181,-16'd6391,-16'd11940,-16'd4427,16'd4633,-16'd7035,-16'd3514,16'd8346,-16'd5199,16'd2387,16'd7986,16'd3713,-16'd7490,16'd1610,-16'd10033,-16'd6106,16'd7532,-16'd4577,-16'd4289,-16'd576,16'd6675,-16'd3091,16'd2704,16'd3078,16'd2881};
dout[92]={ -16'd5271,-16'd7346,16'd6449,16'd5447,16'd4546,16'd5282,-16'd3191,16'd5656,16'd433,-16'd8270,16'd4800,-16'd2408,16'd3719,-16'd4126,-16'd1634,16'd73,-16'd3440,16'd2353,16'd862,16'd3817,16'd2455,16'd5107,-16'd6412,-16'd853,-16'd5654,-16'd15412,16'd2196,-16'd97,-16'd10846,16'd2458,-16'd4315,16'd2530,-16'd5258,-16'd11872,-16'd1658,16'd9419};
dout[93]={ -16'd4835,16'd3225,16'd4992,16'd1125,16'd3231,-16'd3883,-16'd5248,16'd742,16'd5764,-16'd628,16'd6475,-16'd4502,16'd6605,16'd1671,16'd500,-16'd5050,-16'd7037,16'd3272,-16'd7254,-16'd2513,16'd2757,-16'd3766,16'd2084,-16'd8069,16'd7605,-16'd10452,-16'd3189,-16'd3502,-16'd4235,16'd6641,-16'd1910,-16'd9412,-16'd464,16'd5919,-16'd1168,16'd8692};
dout[94]={ -16'd5991,-16'd5700,16'd1292,16'd977,16'd7252,-16'd1158,16'd2205,16'd6236,16'd4863,16'd7943,-16'd1736,-16'd3174,16'd2401,-16'd1282,-16'd4094,16'd552,-16'd5066,-16'd297,-16'd8471,16'd27,16'd696,-16'd5847,-16'd9032,-16'd1485,16'd5267,-16'd5868,16'd3764,16'd1657,16'd3513,-16'd1738,16'd429,-16'd3302,-16'd3351,16'd3676,-16'd827,16'd1146};
dout[95]={ -16'd1200,16'd1272,16'd741,-16'd3513,-16'd3705,16'd6727,-16'd1342,-16'd4251,16'd1046,-16'd766,-16'd1362,-16'd2071,16'd3295,16'd4623,-16'd9453,16'd434,16'd4612,16'd2108,16'd6107,16'd1042,16'd2256,16'd2086,-16'd5700,16'd5344,16'd4638,-16'd2101,16'd1490,16'd3896,-16'd3403,16'd8728,-16'd981,16'd3175,16'd3690,16'd555,16'd1138,-16'd1260};
dout[96]={ 16'd1919,-16'd2510,16'd860,-16'd432,16'd3686,16'd6455,16'd6680,-16'd4089,-16'd8174,16'd1060,16'd2296,16'd2763,16'd1960,16'd459,-16'd7322,16'd5584,-16'd1358,-16'd4459,-16'd2234,16'd3823,-16'd213,-16'd2922,16'd302,16'd6345,-16'd6917,-16'd50,16'd2417,-16'd2794,-16'd6001,-16'd813,-16'd7560,16'd313,16'd240,16'd2586,-16'd292,-16'd1538};
dout[97]={ 16'd1761,16'd3778,-16'd7549,-16'd234,16'd1522,16'd7198,-16'd6705,16'd372,-16'd6354,16'd592,16'd6757,-16'd6335,-16'd3050,-16'd4538,16'd2936,-16'd7998,-16'd3102,-16'd5836,-16'd536,16'd5728,-16'd7650,16'd3090,16'd5124,-16'd1473,-16'd3356,16'd3549,-16'd3837,-16'd565,16'd2962,16'd640,16'd4082,16'd5265,-16'd69,-16'd926,16'd4419,-16'd4019};
dout[98]={ 16'd677,-16'd1888,-16'd9533,-16'd6665,16'd2625,16'd2676,16'd2630,-16'd100,16'd1416,16'd3160,16'd3855,-16'd9647,-16'd2354,-16'd7760,-16'd6247,-16'd3440,16'd926,16'd132,-16'd698,-16'd4866,16'd8219,16'd5184,16'd5206,16'd3901,16'd3943,16'd5820,16'd704,16'd865,16'd3081,16'd3024,16'd3664,-16'd1991,16'd4659,16'd2516,16'd2626,16'd873};
dout[99]={ 16'd2045,-16'd7227,-16'd9070,-16'd6551,-16'd5405,16'd319,-16'd5804,16'd3558,-16'd7637,-16'd3234,-16'd6089,-16'd2236,16'd1951,-16'd7024,16'd4426,-16'd2504,-16'd6368,16'd1227,16'd1840,-16'd1196,-16'd4686,16'd1838,-16'd3150,-16'd7378,16'd1592,16'd3612,-16'd8919,-16'd1155,16'd909,16'd89,16'd2193,-16'd6952,16'd5828,-16'd2751,-16'd2714,-16'd6138};
dout[100]={ -16'd4299,16'd2205,-16'd5967,-16'd5811,-16'd1584,-16'd3072,-16'd6595,16'd9082,16'd5427,-16'd7344,-16'd6678,16'd150,-16'd8890,16'd269,-16'd5338,16'd2352,-16'd11438,16'd5845,16'd662,-16'd1777,-16'd2453,16'd9720,-16'd4881,-16'd8717,-16'd2250,-16'd581,16'd2685,-16'd1815,16'd4578,16'd5486,-16'd2261,-16'd6289,-16'd7113,16'd3732,16'd6557,16'd7358};
dout[101]={ -16'd421,16'd2948,-16'd2062,-16'd5001,16'd7087,-16'd8424,-16'd5149,-16'd3157,16'd4083,-16'd5617,-16'd11637,-16'd6083,16'd5723,-16'd8643,-16'd2728,16'd4336,-16'd1304,16'd3440,16'd7768,-16'd1255,-16'd3759,16'd1967,-16'd9554,-16'd716,-16'd5117,16'd3265,16'd596,16'd1463,-16'd3833,16'd3218,16'd2446,16'd382,-16'd7279,-16'd9368,16'd3363,-16'd6589};
dout[102]={ 16'd5653,16'd5129,-16'd1619,16'd2386,-16'd2209,-16'd2614,-16'd586,-16'd1736,-16'd5814,16'd6365,16'd3256,-16'd7367,-16'd7025,-16'd3582,16'd60,16'd3180,-16'd9015,-16'd2608,16'd1327,-16'd314,-16'd3370,16'd4208,-16'd1461,-16'd2964,-16'd9178,16'd1719,-16'd641,16'd5138,-16'd2086,16'd6950,16'd1616,16'd4385,-16'd798,-16'd4539,-16'd3774,-16'd2436};
dout[103]={ 16'd3134,-16'd8407,16'd5205,-16'd4336,16'd4206,16'd2917,16'd5712,16'd1068,16'd2764,16'd7728,-16'd1493,-16'd1757,-16'd6236,-16'd8424,-16'd3102,-16'd1664,-16'd2902,16'd2994,-16'd2473,16'd3325,16'd4052,16'd3037,-16'd8928,16'd331,-16'd6880,-16'd7222,16'd2926,-16'd4109,-16'd7958,16'd1409,-16'd8070,-16'd2716,16'd4419,16'd4498,-16'd4278,16'd9293};
dout[104]={ 16'd6316,-16'd3541,-16'd8726,-16'd6742,16'd7299,16'd10480,16'd2369,16'd7540,-16'd5094,16'd7978,-16'd6902,16'd3916,-16'd5954,-16'd6512,-16'd2768,16'd2324,16'd7605,16'd5348,16'd3737,-16'd2303,16'd5776,16'd1621,-16'd4055,-16'd4564,16'd5880,16'd6298,16'd7554,16'd1471,-16'd1151,-16'd2381,-16'd9668,-16'd2879,16'd6466,-16'd855,-16'd1743,-16'd389};
dout[105]={ 16'd1918,16'd4159,-16'd6390,-16'd6280,-16'd828,16'd3598,-16'd1230,-16'd3447,16'd1704,16'd726,16'd3967,-16'd2998,-16'd5300,16'd187,16'd843,16'd4772,-16'd961,16'd1921,16'd3636,16'd4707,-16'd1803,16'd5332,16'd3556,-16'd2087,-16'd194,16'd6052,-16'd3346,16'd7533,16'd4469,16'd1633,-16'd8812,-16'd6718,16'd3649,-16'd2802,-16'd2124,-16'd181};
dout[106]={ -16'd4703,-16'd827,-16'd10814,16'd1763,16'd1607,-16'd4575,-16'd4418,16'd2425,-16'd2636,16'd6380,-16'd4740,16'd2802,16'd4562,-16'd2307,16'd83,-16'd4030,16'd5508,-16'd3932,16'd1753,-16'd856,-16'd1163,-16'd3395,16'd4499,16'd2489,16'd5020,-16'd4792,-16'd5611,-16'd6040,16'd3957,16'd4029,-16'd7878,16'd1189,-16'd6119,-16'd2279,-16'd6495,-16'd748};
dout[107]={ -16'd8531,-16'd1651,-16'd1742,-16'd8028,-16'd1556,16'd275,16'd3349,16'd2398,-16'd6961,16'd7281,-16'd6502,-16'd4691,-16'd6375,-16'd1457,16'd3366,-16'd4994,-16'd2451,16'd4310,-16'd5959,16'd2612,-16'd4401,16'd778,16'd5679,-16'd907,-16'd7549,16'd6167,-16'd3375,-16'd2967,16'd2339,-16'd1932,-16'd7229,-16'd7092,-16'd1595,-16'd1472,-16'd2413,16'd6836};
dout[108]={ -16'd1421,-16'd1729,-16'd5896,-16'd6112,16'd5065,-16'd3208,-16'd2161,-16'd6013,16'd5367,16'd2016,16'd4514,16'd8086,16'd3959,16'd6239,-16'd4389,-16'd3808,16'd3310,16'd1439,-16'd8707,-16'd3089,-16'd8236,16'd7167,16'd6333,-16'd10,16'd1890,16'd6813,-16'd5126,-16'd8262,16'd3558,-16'd3048,-16'd4751,-16'd7051,16'd6014,16'd5561,16'd638,-16'd7830};
dout[109]={ 16'd6431,-16'd7302,16'd1495,-16'd1852,16'd2756,-16'd8108,-16'd7785,16'd413,16'd3296,-16'd2819,-16'd2304,16'd6007,16'd1814,-16'd5006,16'd680,16'd8050,16'd1571,16'd6485,16'd4334,16'd5052,-16'd6948,-16'd825,-16'd5995,16'd6745,-16'd4644,-16'd5654,-16'd249,-16'd5556,-16'd2401,-16'd6965,16'd1561,-16'd3544,16'd913,-16'd6508,-16'd4498,16'd2000};
dout[110]={ -16'd6372,-16'd2342,16'd1009,-16'd7061,16'd6435,16'd3176,16'd3323,16'd9312,-16'd3324,16'd189,-16'd17188,16'd8077,16'd4721,16'd97,-16'd7627,16'd6697,-16'd6207,-16'd2658,16'd3824,-16'd1774,-16'd1866,-16'd20,-16'd6485,-16'd3022,-16'd993,-16'd3364,16'd2641,-16'd4468,-16'd6007,16'd9024,-16'd5941,-16'd5162,16'd2533,16'd8660,-16'd4132,16'd8526};
dout[111]={ 16'd4083,16'd989,16'd1044,-16'd394,-16'd37,16'd4030,16'd3202,-16'd3946,-16'd175,16'd5683,-16'd3480,16'd4727,-16'd1838,-16'd12758,16'd2734,16'd279,-16'd2543,-16'd879,16'd2801,16'd888,-16'd2781,16'd9895,-16'd545,-16'd5887,16'd4357,16'd2791,-16'd3282,-16'd1982,16'd1475,-16'd3203,-16'd3964,-16'd3496,-16'd2949,-16'd4336,16'd1404,16'd6335};
dout[112]={ 16'd6682,16'd6033,16'd4722,-16'd2679,16'd43,16'd2401,16'd2704,-16'd2885,-16'd2764,16'd2245,-16'd3879,-16'd8097,-16'd4869,-16'd10431,-16'd1784,-16'd4876,-16'd5234,-16'd5020,-16'd4708,16'd3347,-16'd456,16'd7854,-16'd5799,16'd733,16'd3966,-16'd1534,-16'd4152,-16'd5088,-16'd11887,16'd8401,-16'd3516,16'd2801,-16'd10055,-16'd7700,-16'd10340,16'd547};
dout[113]={ -16'd1498,16'd5340,16'd4492,-16'd5123,16'd9191,16'd3306,-16'd5423,16'd1192,-16'd3178,16'd4203,16'd6827,-16'd4404,16'd4897,16'd3399,16'd494,-16'd3337,-16'd817,16'd1589,-16'd1724,-16'd4329,-16'd2255,16'd2645,16'd2615,-16'd7969,16'd7028,-16'd6747,16'd2688,16'd193,-16'd352,-16'd4252,-16'd6146,16'd5078,16'd3326,16'd1211,16'd1275,-16'd3257};
dout[114]={ 16'd5725,16'd5026,-16'd9832,-16'd6832,16'd779,16'd8503,-16'd1386,-16'd6137,16'd5239,16'd1353,16'd1167,16'd4499,16'd4361,-16'd3567,-16'd7019,-16'd7627,-16'd1467,16'd9,-16'd7011,16'd3113,16'd2264,-16'd1658,-16'd4172,16'd3169,-16'd1830,-16'd1331,16'd9534,16'd3197,16'd1170,16'd10,16'd451,-16'd7661,-16'd2002,-16'd2266,16'd778,-16'd2853};
dout[115]={ 16'd2437,-16'd1780,-16'd10388,-16'd8382,16'd4336,16'd1714,16'd771,16'd7101,-16'd4579,16'd6976,-16'd7590,16'd432,16'd5036,16'd3128,-16'd439,16'd5187,16'd4298,-16'd2563,16'd2807,16'd2737,-16'd4804,16'd1972,16'd4124,-16'd4373,-16'd681,-16'd8185,-16'd3992,-16'd7477,16'd4896,-16'd2925,16'd587,-16'd7141,-16'd5383,-16'd5755,16'd6828,-16'd3643};
dout[116]={ -16'd4018,16'd1347,-16'd8379,-16'd5796,-16'd4487,16'd4783,16'd1220,-16'd4791,16'd4928,-16'd3921,16'd565,-16'd2674,16'd6194,16'd5664,16'd2513,-16'd4959,-16'd776,16'd7310,16'd2817,-16'd7693,-16'd1432,16'd3265,-16'd2903,-16'd2231,16'd2821,16'd872,-16'd5863,-16'd7067,16'd2177,16'd1786,-16'd4025,16'd2928,16'd1191,16'd3397,-16'd6768,16'd2559};
dout[117]={ -16'd1663,16'd89,-16'd6343,16'd772,16'd5077,16'd363,-16'd5860,16'd3200,16'd2881,-16'd367,16'd1647,16'd6177,16'd1501,16'd1184,-16'd8649,16'd3791,-16'd4226,-16'd3473,-16'd3151,16'd2776,-16'd7055,16'd4152,16'd528,-16'd3595,16'd3440,16'd5990,-16'd8030,16'd3000,-16'd4786,-16'd5849,16'd6228,-16'd4817,16'd938,16'd3309,16'd4511,-16'd3797};
dout[118]={ -16'd962,16'd1489,-16'd7682,16'd3322,-16'd1107,16'd1038,-16'd1116,-16'd3162,-16'd3116,16'd1138,-16'd971,16'd4745,16'd7177,16'd5526,-16'd3973,16'd1611,-16'd1852,16'd999,16'd4310,16'd1688,-16'd6657,16'd6227,-16'd7634,16'd4550,16'd809,-16'd5504,-16'd1731,16'd3851,16'd3016,16'd5700,-16'd4481,-16'd345,-16'd666,-16'd7968,16'd1690,-16'd8554};
dout[119]={ -16'd4513,-16'd2631,-16'd1583,16'd2117,16'd2481,-16'd5125,-16'd2056,-16'd6455,-16'd5161,16'd5956,-16'd5405,-16'd2276,16'd5931,-16'd2867,16'd4286,16'd5852,16'd5970,16'd3910,16'd2035,16'd717,16'd8007,-16'd2892,-16'd3884,-16'd6456,-16'd10235,-16'd110,-16'd4691,16'd1815,-16'd2209,-16'd2746,16'd2605,16'd1163,16'd2484,16'd4693,-16'd7081,-16'd73};
dout[120]={ 16'd254,16'd4659,16'd4048,16'd2180,16'd5362,-16'd2680,16'd12281,16'd4106,-16'd7940,16'd817,-16'd11567,-16'd1115,16'd338,-16'd2976,-16'd3221,16'd2004,16'd516,-16'd3635,16'd1907,16'd8036,-16'd1467,16'd7096,-16'd5734,-16'd275,-16'd2941,-16'd7031,16'd6845,-16'd9654,16'd4008,16'd4159,-16'd6934,16'd4412,-16'd2428,-16'd5016,16'd781,16'd6014};
dout[121]={ 16'd7187,16'd278,-16'd1088,-16'd4595,-16'd3861,-16'd2593,16'd5987,16'd2355,-16'd2009,-16'd7134,-16'd7167,16'd7415,-16'd3634,-16'd11522,16'd1562,-16'd1389,-16'd8387,-16'd9753,-16'd4475,16'd5131,16'd3665,16'd568,-16'd6662,-16'd3719,16'd1695,-16'd4394,-16'd1837,-16'd6202,-16'd10465,-16'd5027,-16'd3996,16'd4342,16'd5367,16'd3329,16'd7502,16'd4045};
dout[122]={ 16'd6246,-16'd1827,16'd4277,16'd4389,16'd6666,-16'd1307,16'd4358,-16'd8003,-16'd6488,16'd3934,16'd6483,16'd4388,-16'd8195,-16'd166,-16'd4643,-16'd2906,-16'd4427,-16'd175,16'd997,16'd4035,16'd1165,-16'd27,16'd2910,-16'd5247,-16'd343,-16'd4335,16'd4366,16'd1493,-16'd6762,-16'd3091,-16'd1064,-16'd598,-16'd7799,-16'd4978,16'd2445,16'd4674};
dout[123]={ -16'd703,-16'd4351,16'd7529,-16'd3255,-16'd3903,-16'd1739,16'd1516,16'd5454,-16'd2351,16'd6960,16'd10763,-16'd6137,-16'd1818,-16'd4002,16'd5450,-16'd4019,16'd3757,-16'd5089,16'd5611,16'd506,16'd2185,-16'd3851,16'd4484,-16'd1251,16'd4256,-16'd269,-16'd4545,-16'd6071,16'd4453,-16'd4001,16'd2565,16'd5885,-16'd3593,-16'd1083,16'd1332,-16'd246};
dout[124]={ 16'd4350,16'd7802,16'd5139,-16'd6597,16'd2287,16'd5407,16'd5913,-16'd3314,16'd3785,-16'd4289,16'd6758,-16'd638,16'd3072,16'd2297,-16'd1135,16'd4325,16'd10300,16'd768,16'd1179,-16'd7400,16'd3188,16'd4808,-16'd5800,-16'd6923,16'd4273,-16'd5701,-16'd1517,-16'd1354,16'd4674,-16'd6515,-16'd3278,-16'd3979,-16'd6832,16'd8165,16'd5191,-16'd2825};
dout[125]={ -16'd4482,-16'd4605,16'd3837,-16'd3391,16'd5421,-16'd1525,16'd4645,16'd4939,16'd2832,-16'd4218,16'd987,-16'd4144,16'd2133,-16'd3506,16'd2487,-16'd4177,-16'd4020,-16'd5082,16'd5930,-16'd3640,-16'd2165,-16'd236,-16'd7081,16'd3835,16'd1628,-16'd5558,16'd4551,-16'd1958,16'd5340,16'd2044,16'd2799,-16'd2744,-16'd2734,-16'd2676,16'd1900,-16'd3127};
dout[126]={ -16'd3528,-16'd2261,16'd4748,-16'd8226,16'd3128,-16'd3457,16'd8756,16'd5866,16'd4233,-16'd1321,16'd139,-16'd27,-16'd4979,16'd2359,16'd1383,-16'd6805,16'd4403,16'd36,-16'd6598,-16'd2283,-16'd4073,16'd6925,16'd3308,-16'd3838,-16'd2325,16'd5303,-16'd1344,-16'd5583,-16'd2593,-16'd7855,-16'd3975,16'd3141,-16'd588,-16'd3799,-16'd9408,16'd6092};
dout[127]={ 16'd4243,-16'd1562,-16'd8548,-16'd150,16'd177,-16'd4934,-16'd5945,16'd3047,16'd1248,-16'd1134,-16'd2959,-16'd2549,-16'd602,-16'd4219,16'd2580,-16'd1161,-16'd1861,-16'd1505,-16'd6850,16'd2431,-16'd2265,-16'd961,-16'd2258,16'd3551,-16'd1763,-16'd399,-16'd8183,-16'd7451,-16'd3294,16'd4143,-16'd1471,-16'd5615,-16'd6610,16'd367,16'd2209,-16'd2493};
dout[128]={ -16'd226,-16'd4265,-16'd1937,-16'd5894,16'd3293,-16'd10305,16'd4206,-16'd3581,16'd2648,16'd4780,16'd3073,-16'd5065,-16'd7387,16'd3892,-16'd7757,-16'd3222,16'd1580,16'd4090,16'd3877,-16'd4465,16'd2719,16'd6805,-16'd315,16'd3594,16'd3965,16'd6890,-16'd189,-16'd7520,16'd5896,-16'd3543,-16'd7784,-16'd6080,16'd3365,16'd7298,16'd814,-16'd7237};
dout[129]={ -16'd558,-16'd46,-16'd625,-16'd670,-16'd3226,-16'd3996,16'd3110,-16'd2420,-16'd8073,-16'd2901,16'd2519,16'd4012,-16'd642,16'd1004,-16'd4813,16'd4461,-16'd3397,-16'd4210,-16'd1499,-16'd5126,16'd3827,16'd3603,-16'd1642,16'd3549,-16'd8301,-16'd1301,16'd2928,-16'd1196,16'd6673,-16'd6006,16'd6128,16'd4291,16'd4118,-16'd5223,16'd146,-16'd493};
dout[130]={ -16'd2913,-16'd4524,16'd7067,16'd2310,16'd2875,-16'd3751,16'd10532,16'd10385,16'd6116,16'd7623,-16'd13524,-16'd4199,-16'd9957,-16'd7306,-16'd6931,16'd1682,16'd2878,-16'd4653,-16'd4138,-16'd1361,-16'd4111,-16'd3711,-16'd1518,-16'd8899,-16'd4116,16'd3300,16'd188,16'd2150,-16'd1734,-16'd158,16'd640,16'd1420,-16'd828,-16'd1657,-16'd5933,16'd4228};
dout[131]={ 16'd4683,-16'd1660,-16'd3302,-16'd1832,16'd891,16'd2597,16'd5477,-16'd10238,-16'd7097,-16'd3045,16'd3988,16'd7825,-16'd7750,-16'd1148,16'd4135,16'd1563,-16'd3445,-16'd4203,16'd2250,-16'd6594,16'd5561,16'd430,16'd723,16'd2043,16'd7109,-16'd8008,-16'd2363,-16'd9693,16'd3227,-16'd9483,16'd3786,-16'd962,16'd306,-16'd1740,-16'd4274,16'd109};
dout[132]={ -16'd787,-16'd2637,16'd558,16'd7456,16'd4302,-16'd6008,-16'd875,16'd2800,-16'd3899,16'd8935,16'd2251,16'd6507,-16'd7435,-16'd4846,-16'd285,-16'd8160,16'd2793,-16'd3451,16'd8252,16'd7484,-16'd2753,-16'd4828,16'd1425,-16'd3499,16'd7188,16'd3548,16'd1868,-16'd7413,-16'd3861,-16'd3407,16'd3323,-16'd1062,16'd5602,-16'd8988,-16'd3419,-16'd2009};
dout[133]={ 16'd6124,16'd6900,16'd1972,16'd885,-16'd3872,-16'd601,16'd2768,-16'd4503,-16'd2851,-16'd948,16'd3501,16'd3863,-16'd6869,-16'd10413,16'd1006,16'd2921,16'd2763,-16'd7455,-16'd3951,16'd5539,16'd3349,16'd5613,16'd4659,-16'd7475,16'd1301,-16'd4803,-16'd4345,-16'd7186,-16'd4412,-16'd5486,-16'd1328,-16'd329,-16'd4159,16'd3512,16'd6039,-16'd3403};
dout[134]={ 16'd4263,16'd2947,-16'd1741,16'd4971,-16'd2822,16'd1784,-16'd3003,16'd3966,-16'd3124,16'd4439,-16'd6791,16'd0,-16'd5889,16'd1025,16'd2697,16'd5888,-16'd2660,16'd3159,-16'd7172,-16'd2125,16'd4974,16'd4324,16'd2132,16'd483,-16'd1513,-16'd4227,-16'd2994,-16'd3931,-16'd1203,-16'd5156,-16'd7681,16'd2126,-16'd3063,-16'd820,-16'd3018,-16'd11536};
dout[135]={ -16'd2597,16'd1253,-16'd2098,-16'd5979,-16'd9059,-16'd2251,-16'd1495,-16'd5935,16'd3897,16'd4948,16'd3909,16'd1116,-16'd3668,-16'd7853,16'd761,-16'd2245,-16'd3391,-16'd6640,16'd6309,16'd2777,-16'd1691,-16'd53,-16'd3193,16'd3802,16'd5357,-16'd3515,16'd4643,16'd1870,16'd3839,-16'd2700,16'd1710,16'd4296,-16'd3632,16'd7893,16'd528,16'd6456};
dout[136]={ 16'd4168,-16'd1905,16'd1256,-16'd988,16'd2994,16'd2091,-16'd5861,16'd4927,-16'd6129,-16'd2502,16'd556,-16'd936,-16'd5178,16'd5368,-16'd8858,-16'd5359,-16'd3280,-16'd5640,-16'd3121,16'd502,16'd1775,16'd5442,16'd7123,-16'd3293,-16'd1948,16'd4679,16'd2718,16'd1764,-16'd1645,-16'd5659,16'd1592,16'd499,16'd5187,-16'd4315,-16'd1086,-16'd5420};
dout[137]={ 16'd1715,-16'd2602,-16'd2514,16'd1382,16'd1258,-16'd1991,16'd5794,-16'd1392,-16'd5080,16'd2713,16'd538,-16'd134,-16'd4704,16'd5935,16'd5229,-16'd1112,-16'd1108,-16'd729,16'd5150,-16'd5714,-16'd8082,-16'd842,16'd7384,16'd2794,16'd2832,16'd5713,-16'd7215,16'd3490,16'd5446,16'd5217,16'd6096,16'd2626,16'd571,-16'd1933,16'd880,-16'd7625};
dout[138]={ -16'd5557,-16'd3955,16'd1601,-16'd3121,-16'd5394,-16'd5048,16'd3576,-16'd2446,-16'd3937,16'd832,-16'd248,-16'd2485,-16'd7106,-16'd1950,-16'd7268,16'd5793,-16'd1042,16'd6056,16'd2450,16'd2347,-16'd8474,-16'd947,16'd5820,-16'd4600,16'd4097,16'd10192,16'd3890,-16'd276,-16'd4848,16'd2375,-16'd6497,16'd3625,-16'd5787,-16'd4778,16'd4722,-16'd4823};
dout[139]={ -16'd6132,16'd1878,-16'd1546,-16'd2137,-16'd3693,16'd3793,16'd1159,-16'd1353,16'd3212,16'd1006,16'd1585,16'd4001,-16'd1954,16'd5069,-16'd2526,-16'd5478,16'd600,16'd2064,16'd2401,16'd2897,-16'd4053,-16'd3576,16'd4720,-16'd3034,16'd7412,-16'd1280,-16'd4529,-16'd2874,16'd2078,-16'd2957,16'd259,16'd2204,16'd166,-16'd3616,-16'd7723,-16'd5710};
dout[140]={ -16'd4808,16'd5362,-16'd2018,-16'd5178,-16'd3930,-16'd8673,-16'd2279,16'd8052,-16'd7186,16'd8415,16'd4172,-16'd6419,-16'd13589,-16'd10342,16'd5442,16'd6546,16'd6021,-16'd1921,16'd6247,16'd5461,16'd907,16'd6511,16'd1660,-16'd1396,-16'd70,16'd3845,16'd3565,-16'd7382,16'd5570,-16'd9009,-16'd5442,16'd99,16'd5445,-16'd4954,16'd5286,16'd10578};
dout[141]={ -16'd2535,-16'd5594,16'd6044,16'd2812,-16'd3677,-16'd6487,-16'd2609,-16'd8417,16'd4740,16'd2472,16'd8020,-16'd2974,16'd2176,-16'd5645,16'd1300,16'd3269,-16'd2093,16'd4458,16'd8120,-16'd3895,16'd6508,16'd3634,16'd5345,-16'd2797,-16'd2427,-16'd6388,16'd338,-16'd538,-16'd6513,-16'd4648,-16'd777,-16'd1429,-16'd1442,-16'd3367,-16'd5106,16'd646};
dout[142]={ 16'd313,-16'd2016,-16'd2927,16'd7690,-16'd6101,16'd635,-16'd5407,-16'd1181,-16'd2946,-16'd2019,-16'd159,16'd2327,-16'd2303,-16'd5619,16'd3581,16'd3570,16'd5487,16'd6198,16'd8204,-16'd3695,16'd1382,-16'd7271,-16'd5778,-16'd8637,16'd2617,-16'd7145,16'd1476,16'd1264,-16'd9091,-16'd6908,-16'd2658,16'd1805,16'd4517,-16'd9142,16'd4908,16'd1651};
dout[143]={ 16'd6065,16'd3422,-16'd2055,-16'd1940,-16'd3271,16'd3921,-16'd7851,16'd9032,-16'd28,16'd2776,16'd4962,16'd8974,16'd4732,-16'd1768,16'd5581,-16'd6125,16'd4732,16'd829,16'd4095,16'd4104,16'd1621,16'd2715,-16'd4983,-16'd9877,16'd580,16'd1195,16'd6585,-16'd10308,-16'd3983,-16'd4795,16'd1913,-16'd5906,-16'd3937,-16'd1379,16'd8457,-16'd9432};
dout[144]={ 16'd4894,16'd1740,-16'd158,16'd5460,-16'd3230,-16'd3622,-16'd3996,-16'd866,16'd2199,16'd6645,-16'd4364,-16'd4787,-16'd3366,16'd392,-16'd1852,16'd4255,16'd2293,16'd394,-16'd7730,-16'd1716,-16'd4305,16'd1284,-16'd2868,16'd136,-16'd8695,-16'd5258,-16'd3357,-16'd3678,16'd4680,-16'd5858,-16'd8022,-16'd5887,-16'd6384,16'd479,-16'd1304,16'd1221};
dout[145]={ -16'd543,16'd5498,-16'd1285,-16'd7276,-16'd4038,16'd2143,16'd1586,16'd4112,-16'd980,16'd8083,16'd6301,16'd8846,-16'd1780,-16'd8216,16'd3392,16'd3015,-16'd422,-16'd843,-16'd3659,-16'd464,-16'd3717,-16'd2591,-16'd3149,16'd5762,-16'd7293,-16'd4416,-16'd7622,16'd3204,16'd2866,-16'd9355,-16'd3037,-16'd325,16'd1083,16'd3015,16'd2680,-16'd7157};
dout[146]={ -16'd2873,-16'd2114,-16'd1248,-16'd7116,-16'd645,16'd3157,-16'd7545,-16'd1315,-16'd5895,16'd2571,16'd1939,-16'd6098,-16'd3450,-16'd8770,-16'd3534,-16'd1547,-16'd5024,-16'd6670,-16'd3294,16'd1981,-16'd10408,-16'd3699,-16'd4535,-16'd1132,-16'd623,-16'd7225,16'd1463,-16'd6078,-16'd4082,16'd2016,-16'd910,-16'd2746,-16'd6893,16'd394,-16'd7246,-16'd1324};
dout[147]={ -16'd5031,16'd6121,16'd2449,16'd6514,16'd3066,-16'd8050,16'd4909,-16'd6393,16'd1647,-16'd4721,16'd7962,16'd6790,16'd532,16'd2107,-16'd1062,-16'd6182,16'd210,16'd3912,16'd4337,16'd5380,-16'd6992,16'd2651,16'd6948,16'd4598,16'd1713,16'd4001,-16'd3515,16'd2113,16'd1181,-16'd5582,16'd6196,-16'd6206,16'd686,-16'd4062,-16'd448,16'd1945};
dout[148]={ 16'd3501,16'd2473,16'd1735,-16'd6105,16'd1653,-16'd2839,-16'd9163,16'd708,-16'd6779,-16'd1806,-16'd2349,-16'd5268,16'd5355,-16'd5066,16'd3721,-16'd4228,16'd1101,16'd5400,-16'd4483,16'd5213,16'd1659,16'd2680,16'd1711,16'd5930,-16'd837,-16'd3580,16'd2770,16'd1265,-16'd3879,-16'd394,16'd5743,16'd1572,-16'd1668,-16'd154,-16'd5612,-16'd8716};
dout[149]={ -16'd2033,16'd4853,-16'd5445,-16'd534,-16'd2377,16'd5930,16'd5709,16'd5180,16'd6191,16'd3363,-16'd3860,-16'd6051,16'd6105,16'd3963,-16'd3584,-16'd890,16'd4782,-16'd3708,-16'd3569,16'd1929,-16'd5566,16'd7771,16'd5162,16'd3903,-16'd1259,16'd8822,-16'd4664,-16'd2594,16'd3617,-16'd3688,16'd1833,-16'd6359,-16'd4528,16'd5339,-16'd3300,-16'd7453};
dout[150]={ -16'd4054,-16'd3960,16'd6302,16'd5262,-16'd3213,16'd175,-16'd7831,16'd4096,-16'd1379,16'd3138,16'd242,16'd935,-16'd6060,-16'd7647,-16'd1680,-16'd2051,-16'd788,16'd6671,16'd2047,-16'd1815,-16'd1760,16'd1450,16'd4215,-16'd198,16'd314,-16'd959,-16'd464,16'd385,16'd3650,-16'd15219,-16'd8764,16'd1652,16'd758,-16'd34,16'd8000,16'd1661};
dout[151]={ -16'd4117,-16'd480,-16'd6486,16'd4874,16'd2806,16'd623,16'd4434,16'd28,-16'd3276,16'd145,16'd3439,16'd777,16'd5860,16'd536,-16'd3906,-16'd3026,-16'd2217,-16'd4381,16'd7289,16'd3068,16'd830,16'd3736,16'd3559,-16'd9794,16'd5065,16'd4210,-16'd4886,-16'd6086,-16'd408,-16'd4670,16'd4541,-16'd395,16'd6411,-16'd2095,-16'd3726,16'd6039};
dout[152]={ 16'd5046,16'd2241,16'd4162,16'd11583,16'd2870,-16'd1029,-16'd9475,16'd1450,16'd1845,16'd11251,16'd6668,16'd2882,-16'd6987,16'd3100,-16'd3028,16'd2681,-16'd476,-16'd5904,16'd6667,16'd812,-16'd2862,16'd1151,16'd493,-16'd5101,-16'd1578,-16'd10436,16'd2037,16'd55,-16'd6720,-16'd5490,16'd522,16'd1078,16'd8228,16'd5360,16'd795,-16'd3346};
dout[153]={ 16'd4942,-16'd7023,16'd3403,16'd9148,-16'd5557,16'd4287,-16'd7175,16'd9284,-16'd7538,16'd8008,16'd5723,-16'd5272,16'd6581,-16'd5090,-16'd668,-16'd7845,-16'd3952,16'd2121,16'd639,16'd6029,16'd2173,16'd5454,-16'd1603,-16'd3923,16'd3379,-16'd2615,16'd4149,16'd260,-16'd2893,16'd782,-16'd8614,16'd4761,16'd5560,-16'd4451,16'd2403,-16'd7503};
dout[154]={ 16'd1273,-16'd681,16'd4294,-16'd5122,16'd320,-16'd830,-16'd10712,-16'd6193,16'd4658,-16'd9244,-16'd6898,16'd1758,16'd925,-16'd6947,-16'd2117,-16'd1965,-16'd3812,-16'd1716,16'd1968,16'd6232,16'd6243,-16'd2867,16'd1489,16'd4628,16'd2236,-16'd6178,-16'd264,16'd658,-16'd312,-16'd6416,16'd488,-16'd4383,-16'd386,-16'd818,16'd2882,16'd683};
dout[155]={ -16'd1742,16'd5041,16'd5883,-16'd567,16'd294,-16'd6003,-16'd1603,-16'd3671,-16'd3834,-16'd6887,-16'd5133,-16'd2335,-16'd5219,-16'd7115,-16'd2169,16'd4341,-16'd97,-16'd2669,-16'd6291,16'd959,16'd3143,16'd1978,16'd2558,16'd106,16'd1834,-16'd6760,16'd5304,16'd7004,16'd5822,-16'd3623,-16'd1289,16'd4351,-16'd293,-16'd352,-16'd615,16'd384};
dout[156]={ -16'd7280,16'd351,16'd4314,-16'd7916,-16'd7429,16'd4744,16'd629,-16'd3493,-16'd651,-16'd3866,-16'd4180,16'd6141,16'd4271,-16'd2110,16'd741,-16'd6418,-16'd4118,-16'd4929,16'd6891,16'd1168,16'd4419,16'd189,-16'd4965,16'd4287,16'd4116,16'd4478,-16'd7173,16'd3442,-16'd221,16'd5009,-16'd4125,-16'd7806,16'd1789,16'd5094,-16'd3945,-16'd4752};
dout[157]={ -16'd8918,16'd3849,-16'd1808,16'd907,-16'd2278,-16'd5504,-16'd5066,-16'd3729,16'd4711,16'd5151,-16'd2942,-16'd3260,16'd4359,16'd4936,-16'd4140,16'd3780,-16'd2708,-16'd5743,16'd2640,16'd6330,-16'd255,16'd5894,-16'd4097,16'd6100,16'd3299,-16'd4187,-16'd181,16'd7034,-16'd3912,-16'd1047,16'd2102,-16'd2471,16'd7859,16'd4099,16'd1441,-16'd541};
dout[158]={ -16'd6499,-16'd4306,16'd408,16'd7369,16'd575,16'd6925,-16'd8243,-16'd2653,-16'd1218,-16'd4482,16'd3833,16'd1266,-16'd758,16'd384,16'd6134,16'd5392,-16'd7198,-16'd7402,-16'd1592,16'd4715,-16'd9171,16'd2421,16'd147,-16'd5848,16'd5857,16'd1063,16'd4949,16'd2173,16'd5789,16'd2720,16'd3947,-16'd7617,-16'd1010,-16'd2351,-16'd4909,-16'd2423};
dout[159]={ -16'd1243,16'd3293,-16'd2177,16'd4635,16'd7059,-16'd2852,16'd804,-16'd5609,16'd368,-16'd5481,-16'd5,16'd1227,16'd3456,16'd5391,-16'd2931,-16'd6286,16'd1829,-16'd2379,16'd1641,16'd2035,-16'd1436,16'd33,16'd1923,16'd4244,16'd7360,16'd7119,16'd2886,-16'd4021,-16'd5041,16'd2207,-16'd3583,-16'd4795,-16'd1674,16'd2417,-16'd1644,-16'd5472};
dout[160]={ 16'd4676,16'd3218,-16'd5419,16'd4368,16'd5057,16'd2347,-16'd9508,16'd1199,-16'd3788,-16'd1144,-16'd3191,16'd2139,-16'd10528,-16'd9882,16'd7479,16'd5567,16'd5625,16'd6393,16'd369,-16'd1063,-16'd6708,16'd142,-16'd6794,-16'd5050,16'd3097,16'd6042,-16'd5514,16'd3015,16'd4279,-16'd10644,-16'd2166,-16'd3553,16'd3891,-16'd2943,16'd706,-16'd1115};
dout[161]={ 16'd161,16'd5119,16'd1960,16'd6116,-16'd8346,-16'd396,16'd396,16'd8910,16'd207,16'd6705,-16'd8755,-16'd4658,-16'd3468,-16'd10340,-16'd7013,16'd6192,-16'd3330,16'd4632,16'd2684,16'd6350,-16'd2120,-16'd5650,-16'd5116,-16'd11842,-16'd1411,-16'd4471,16'd838,-16'd3343,16'd3352,-16'd6110,-16'd2419,-16'd2398,-16'd4607,-16'd6723,-16'd3505,-16'd3072};
dout[162]={ 16'd3340,-16'd9389,-16'd10486,16'd6241,16'd329,-16'd4502,-16'd4856,16'd9000,-16'd1381,16'd4789,-16'd7410,16'd5261,-16'd2096,16'd421,-16'd1338,-16'd3078,-16'd5558,16'd7688,16'd3292,16'd3640,-16'd5663,-16'd10660,16'd2124,-16'd637,16'd1704,-16'd5497,16'd4921,16'd5673,-16'd3158,16'd4523,-16'd6979,16'd2588,-16'd2859,16'd6172,16'd8338,16'd5057};
dout[163]={ -16'd3841,-16'd8609,-16'd7355,16'd6873,16'd2250,-16'd5734,16'd1181,16'd5173,-16'd5453,-16'd7061,-16'd1226,-16'd4057,16'd3680,-16'd10553,-16'd1476,-16'd2469,16'd2373,-16'd643,16'd6448,16'd6136,-16'd810,-16'd4954,16'd4841,-16'd381,-16'd5979,16'd880,-16'd3305,16'd4533,16'd7701,-16'd1040,16'd4069,-16'd2813,-16'd3357,-16'd6045,16'd5753,-16'd985};
dout[164]={ 16'd118,16'd4039,16'd2902,-16'd1006,-16'd5462,16'd1364,-16'd6078,-16'd5138,16'd1507,-16'd11383,16'd932,16'd1823,16'd5388,-16'd8618,16'd7534,-16'd6798,16'd7499,16'd4197,16'd3552,16'd3178,-16'd305,-16'd5439,-16'd1945,-16'd2678,-16'd5202,-16'd2943,-16'd8,16'd7441,16'd2975,16'd2212,-16'd10041,-16'd318,16'd775,16'd3885,-16'd3082,-16'd9733};
dout[165]={ 16'd5073,-16'd402,16'd1167,16'd3641,16'd2243,-16'd6430,-16'd3688,16'd3129,-16'd1406,16'd278,16'd3221,16'd4211,-16'd2620,-16'd2979,16'd6378,-16'd1239,-16'd4486,-16'd3109,16'd5253,-16'd2233,-16'd1537,-16'd2268,-16'd118,-16'd856,16'd193,-16'd514,16'd783,16'd3577,16'd5325,16'd4740,-16'd7558,16'd2270,-16'd1026,16'd2828,-16'd3701,-16'd6559};
dout[166]={ 16'd2327,16'd3894,16'd2961,16'd1867,16'd2283,-16'd3299,-16'd794,-16'd4890,16'd3938,16'd6164,16'd4893,-16'd7954,16'd6365,16'd4044,16'd5766,16'd6341,16'd3382,-16'd11388,-16'd1918,16'd717,-16'd4068,-16'd3754,-16'd220,-16'd18,16'd620,-16'd4747,-16'd6894,16'd1076,16'd6849,16'd4466,16'd4153,16'd2617,16'd2277,16'd476,16'd5962,16'd2257};
dout[167]={ 16'd3976,-16'd6793,-16'd7512,16'd3479,16'd487,16'd2575,-16'd3638,-16'd7205,-16'd2789,16'd1970,-16'd2080,-16'd4665,-16'd1457,16'd3702,16'd6432,16'd1923,-16'd3176,-16'd410,-16'd1784,-16'd654,-16'd6464,16'd6266,16'd2967,-16'd1406,16'd2478,16'd3405,-16'd3827,-16'd1211,-16'd3057,-16'd7003,16'd5401,-16'd8787,16'd8988,16'd7076,-16'd5728,-16'd6214};
dout[168]={ -16'd865,-16'd4338,16'd910,-16'd1111,-16'd7015,16'd1171,16'd282,16'd446,16'd584,16'd658,-16'd3938,-16'd1847,16'd3616,-16'd3797,-16'd480,-16'd6168,16'd5237,-16'd6848,-16'd1807,-16'd5058,-16'd8738,-16'd4525,16'd239,16'd3751,16'd2234,-16'd996,-16'd947,-16'd1162,-16'd8294,-16'd4130,-16'd2761,16'd2915,-16'd4737,16'd1093,-16'd1894,-16'd3423};
dout[169]={ 16'd4525,16'd1691,-16'd963,-16'd2294,-16'd3707,-16'd3189,-16'd5763,16'd2810,16'd2346,16'd5333,-16'd6389,16'd4471,-16'd2790,-16'd1114,-16'd4793,-16'd7239,16'd1455,16'd6259,16'd1752,-16'd5773,-16'd6637,-16'd6084,-16'd6429,-16'd1126,-16'd1911,-16'd3595,16'd4147,16'd7565,-16'd2448,-16'd5517,-16'd3716,-16'd7111,16'd923,16'd5308,16'd8150,16'd5288};
dout[170]={ 16'd675,16'd2871,-16'd1070,16'd1072,16'd4258,-16'd6037,16'd678,16'd1163,-16'd3255,16'd4239,-16'd2427,-16'd2593,16'd6915,-16'd1305,-16'd3086,16'd4340,-16'd2129,-16'd5676,-16'd791,-16'd1918,16'd2377,-16'd6028,-16'd6594,16'd5563,16'd4156,-16'd4323,-16'd2351,16'd103,-16'd5421,-16'd7692,-16'd3855,16'd7150,-16'd8427,-16'd2085,16'd6329,16'd4333};
dout[171]={ -16'd1171,16'd396,-16'd4510,16'd4275,16'd1840,16'd5926,-16'd2359,16'd3631,16'd3271,16'd2457,-16'd11176,-16'd31,16'd4629,-16'd3219,-16'd2022,16'd879,16'd4891,16'd5018,16'd298,16'd450,-16'd8273,16'd2412,-16'd627,16'd2,16'd4790,16'd585,-16'd8182,16'd4980,-16'd2627,16'd5912,-16'd992,16'd1789,-16'd2913,-16'd6905,16'd2194,-16'd2729};
dout[172]={ -16'd5570,16'd3547,-16'd1700,-16'd1286,16'd446,16'd4917,16'd3815,-16'd3835,16'd1791,16'd4288,-16'd7595,-16'd4862,16'd6488,-16'd5018,-16'd11190,-16'd6127,16'd370,16'd3649,-16'd4862,-16'd4659,-16'd1133,-16'd8656,16'd5039,-16'd5831,-16'd3308,-16'd1216,16'd4653,16'd3630,-16'd379,16'd1668,-16'd4773,16'd4698,16'd10446,-16'd4602,16'd3660,-16'd2985};
dout[173]={ 16'd4452,-16'd8567,-16'd6492,16'd309,-16'd4421,16'd4324,16'd3240,16'd5734,16'd2436,-16'd2615,16'd5875,16'd2843,16'd303,-16'd2207,-16'd2909,16'd4709,16'd2643,-16'd4572,16'd2640,-16'd568,-16'd84,-16'd6336,16'd1725,-16'd2309,16'd377,-16'd708,-16'd5053,-16'd3734,-16'd2620,-16'd5356,-16'd8026,16'd4704,16'd4935,-16'd5197,16'd2324,-16'd9607};
dout[174]={ 16'd2727,16'd1315,16'd6155,16'd5690,-16'd1362,-16'd3389,16'd2917,16'd4958,-16'd4069,-16'd4128,-16'd2402,-16'd869,-16'd7301,-16'd4928,16'd5076,-16'd7979,-16'd2926,-16'd887,16'd2869,-16'd4199,16'd7446,-16'd4129,16'd4227,16'd5989,16'd2838,-16'd5871,-16'd5772,16'd5473,16'd773,16'd254,-16'd8204,16'd5556,16'd6713,16'd1934,-16'd4619,16'd2410};
dout[175]={ -16'd3196,-16'd1163,-16'd5230,16'd1115,-16'd2278,-16'd2392,-16'd4999,-16'd727,16'd3270,-16'd4300,-16'd3628,-16'd7031,16'd1489,-16'd857,16'd3133,-16'd5775,16'd871,16'd957,16'd1544,16'd2070,16'd296,-16'd2581,-16'd529,16'd7850,-16'd848,-16'd6590,16'd4812,16'd1220,-16'd4844,-16'd3783,-16'd5947,-16'd8020,-16'd5308,-16'd119,-16'd2531,-16'd10693};
dout[176]={ 16'd5585,16'd3447,16'd5324,-16'd2195,-16'd6569,16'd4439,16'd6720,-16'd2635,16'd1581,16'd3411,-16'd8422,-16'd9276,16'd5236,-16'd6300,16'd2308,-16'd4478,16'd1772,-16'd1257,16'd1052,16'd5838,16'd4679,-16'd3407,16'd7453,16'd5343,-16'd5006,-16'd7665,-16'd6954,16'd4048,16'd6297,16'd743,-16'd3295,-16'd3465,16'd6354,-16'd3054,-16'd4477,-16'd10610};
dout[177]={ -16'd889,-16'd1471,-16'd1291,-16'd2460,-16'd7060,16'd2471,-16'd2025,16'd1633,-16'd6272,-16'd848,-16'd5145,-16'd2055,-16'd5674,-16'd393,-16'd262,16'd4087,-16'd5161,-16'd10927,16'd3936,16'd3992,16'd5470,-16'd1221,16'd4646,-16'd3572,-16'd1867,-16'd1590,16'd1181,-16'd391,16'd1010,-16'd79,16'd2146,16'd1047,-16'd1931,-16'd4244,16'd2689,16'd4057};
dout[178]={ -16'd5423,16'd3943,-16'd6451,16'd5032,16'd5575,-16'd78,-16'd3377,16'd5421,-16'd1889,-16'd396,-16'd1467,-16'd4630,16'd5105,16'd2682,-16'd2929,-16'd4191,16'd4234,16'd974,16'd1818,-16'd5355,16'd1827,16'd2682,-16'd3811,-16'd5497,16'd4973,16'd530,16'd5975,16'd4988,16'd783,-16'd4240,-16'd4113,-16'd6963,-16'd3431,-16'd5324,16'd1481,-16'd5753};
dout[179]={ -16'd8061,-16'd4283,16'd4605,16'd3083,16'd2067,16'd3971,-16'd16,16'd6258,16'd3693,-16'd8482,-16'd3218,-16'd9111,16'd2697,16'd3638,16'd1846,-16'd7988,16'd2454,16'd4289,16'd135,-16'd28,16'd2037,16'd6894,-16'd1415,16'd5280,-16'd777,16'd1854,16'd3532,-16'd7946,-16'd132,-16'd2732,-16'd3172,-16'd6305,-16'd3388,16'd3812,-16'd556,-16'd2290};
dout[180]={ 16'd854,-16'd8349,-16'd7380,16'd4750,-16'd6157,-16'd6340,-16'd4996,-16'd8331,16'd4029,16'd2677,-16'd11815,16'd734,16'd5176,-16'd2097,16'd7162,16'd7207,-16'd1254,16'd910,-16'd5222,-16'd7036,16'd2632,16'd2663,16'd3794,16'd5281,-16'd1728,16'd1818,16'd900,16'd6626,16'd204,-16'd6402,-16'd2441,16'd5206,-16'd929,16'd5071,16'd3433,-16'd160};
dout[181]={ 16'd2904,-16'd7687,16'd5041,-16'd6205,-16'd5466,-16'd7134,-16'd4369,16'd7040,-16'd5170,16'd4191,-16'd2033,16'd2106,16'd3032,-16'd7861,16'd5269,16'd3327,-16'd5790,16'd2944,-16'd6356,-16'd10296,16'd5113,-16'd7534,16'd980,-16'd12689,-16'd1329,-16'd350,-16'd2766,16'd5088,16'd2671,16'd351,16'd5594,-16'd557,-16'd4738,-16'd4903,16'd4525,16'd6637};
dout[182]={ 16'd5459,-16'd619,-16'd2034,16'd5618,-16'd6054,-16'd2301,16'd7087,16'd1916,-16'd2354,16'd1586,-16'd8641,-16'd2503,16'd4696,-16'd4293,-16'd3066,-16'd3766,-16'd3372,16'd2336,-16'd7840,-16'd2377,16'd7591,-16'd1753,-16'd4926,-16'd389,-16'd6101,-16'd4519,-16'd2553,16'd6447,-16'd2379,16'd4298,-16'd1031,16'd4923,16'd588,-16'd1851,16'd3901,-16'd4352};
dout[183]={ -16'd5769,-16'd3736,16'd4831,-16'd1214,-16'd1047,-16'd8863,16'd6113,16'd8415,16'd3878,-16'd5138,16'd4921,-16'd4383,16'd893,16'd1342,-16'd701,-16'd6448,16'd7510,16'd2584,16'd5064,16'd4118,16'd310,16'd4142,-16'd4502,16'd2568,16'd3823,16'd472,16'd3508,-16'd4659,16'd4145,-16'd1360,16'd7687,16'd2312,16'd2043,16'd1047,-16'd5377,-16'd8810};
dout[184]={ 16'd2833,-16'd4089,-16'd4239,16'd3657,-16'd5257,16'd2819,-16'd4591,-16'd1776,16'd5408,-16'd10211,-16'd710,16'd1147,-16'd7534,16'd3394,16'd8763,16'd1595,-16'd3760,-16'd848,16'd3362,16'd2933,16'd7029,16'd5617,16'd2172,16'd1482,-16'd2132,-16'd3151,-16'd9567,-16'd6632,-16'd2190,16'd20,-16'd1110,-16'd3393,-16'd4728,-16'd1730,-16'd4286,-16'd9607};
dout[185]={ -16'd4187,16'd2565,16'd4152,16'd8333,-16'd6169,-16'd3775,16'd4011,-16'd4269,-16'd5460,16'd2977,16'd3475,-16'd2662,16'd4686,16'd4876,16'd3725,16'd561,16'd6763,-16'd3634,-16'd7185,16'd5545,16'd1154,-16'd6114,16'd4446,-16'd2112,16'd4453,-16'd6767,-16'd4522,-16'd548,16'd780,-16'd1249,16'd4697,16'd3597,-16'd4724,16'd1659,-16'd5853,-16'd8532};
dout[186]={ 16'd4783,-16'd2354,-16'd6980,16'd3181,16'd3735,-16'd2957,16'd7118,-16'd1199,16'd3232,16'd839,-16'd4595,16'd2324,16'd244,-16'd2769,16'd5820,-16'd290,-16'd7312,-16'd6931,-16'd713,-16'd6669,16'd5366,16'd3848,-16'd4615,16'd2794,16'd1752,16'd2455,-16'd1614,-16'd8365,-16'd5909,16'd2626,16'd5647,-16'd5648,16'd2726,-16'd2357,16'd5010,-16'd1430};
dout[187]={ -16'd5408,16'd30,16'd1402,16'd5552,16'd2307,16'd1653,16'd4517,16'd2379,-16'd5388,-16'd6082,16'd963,-16'd10398,16'd1390,16'd945,-16'd5196,-16'd5851,16'd4177,16'd127,-16'd152,-16'd7018,-16'd7900,-16'd4512,16'd5087,16'd2787,16'd6726,16'd6118,-16'd4874,-16'd57,16'd2565,-16'd2739,-16'd3566,16'd5903,16'd6293,-16'd1784,16'd3511,-16'd5713};
dout[188]={ -16'd357,-16'd6938,16'd5459,16'd758,-16'd7905,-16'd2721,16'd178,16'd4785,-16'd6353,-16'd8651,16'd2938,-16'd921,-16'd3753,16'd2596,16'd7826,16'd2693,16'd1763,16'd8268,-16'd5573,-16'd290,-16'd5799,16'd4769,-16'd5996,16'd603,16'd2012,-16'd7333,16'd1592,16'd576,-16'd7956,16'd2463,-16'd3467,16'd2931,16'd2550,-16'd8645,16'd3128,-16'd525};
dout[189]={ -16'd6960,-16'd1936,-16'd2292,-16'd1272,16'd3161,16'd7293,-16'd5453,16'd961,16'd2840,16'd1828,-16'd6195,-16'd6251,-16'd1860,-16'd5749,16'd8,16'd3203,16'd6090,16'd763,16'd2695,16'd6671,-16'd8167,16'd5356,16'd1055,-16'd7944,-16'd6679,16'd3859,-16'd3640,16'd3798,16'd483,16'd1083,16'd7679,16'd2236,16'd880,16'd4059,16'd1019,-16'd4223};
dout[190]={ 16'd1964,-16'd8830,-16'd3957,-16'd1737,16'd7803,16'd6208,-16'd3698,16'd1183,-16'd776,16'd5747,-16'd5901,-16'd4153,16'd27,-16'd8450,-16'd529,-16'd7732,-16'd8467,16'd3425,-16'd9605,-16'd4684,16'd3039,-16'd8383,-16'd1888,16'd278,-16'd630,16'd6644,-16'd4516,-16'd6710,16'd1865,16'd424,16'd1860,-16'd5013,16'd1648,16'd7452,16'd1138,-16'd4473};
dout[191]={ 16'd3542,-16'd1458,-16'd6862,-16'd1306,-16'd7160,-16'd8986,-16'd436,16'd4059,16'd7725,-16'd3123,16'd4837,-16'd983,16'd8574,-16'd6806,16'd4894,-16'd2532,-16'd1898,-16'd5194,-16'd2789,-16'd4045,16'd389,-16'd7429,-16'd5164,-16'd3451,16'd112,16'd643,16'd2216,16'd2317,16'd10,16'd3162,16'd192,16'd1468,-16'd4537,-16'd9213,16'd2851,16'd6771};
dout[192]={ 16'd2696,-16'd10845,16'd1088,-16'd2630,16'd2022,-16'd7202,-16'd2782,-16'd331,16'd3444,-16'd6535,16'd2183,16'd276,16'd10065,16'd955,16'd428,16'd4378,-16'd2993,16'd1275,-16'd8474,-16'd9138,-16'd1483,-16'd6775,-16'd574,-16'd163,-16'd2145,16'd1544,-16'd9223,-16'd796,16'd2784,16'd4123,16'd2700,-16'd6193,-16'd909,-16'd2169,-16'd6036,-16'd4220};
dout[193]={ -16'd2522,-16'd9851,-16'd5566,-16'd4333,16'd8019,-16'd3362,16'd1805,16'd583,16'd2179,-16'd12817,16'd189,16'd1433,-16'd4544,-16'd9091,16'd3960,16'd2429,-16'd5056,-16'd6383,16'd3193,-16'd6707,16'd2143,-16'd5360,-16'd7836,-16'd2349,-16'd8816,-16'd4906,-16'd5344,-16'd3392,-16'd2650,16'd5355,16'd2264,-16'd2400,16'd6537,-16'd4224,-16'd9794,16'd4265};
dout[194]={ 16'd6685,16'd5313,-16'd569,-16'd4569,-16'd7619,-16'd72,16'd78,16'd10936,-16'd4802,-16'd4546,-16'd6593,-16'd632,16'd1967,16'd1160,16'd7069,-16'd6586,-16'd3030,16'd7126,16'd9499,16'd9582,-16'd5849,16'd5246,-16'd8822,16'd2579,16'd495,-16'd5227,16'd5169,16'd821,16'd4719,-16'd2048,16'd3614,16'd7366,16'd27,-16'd2156,-16'd8127,16'd4656};
dout[195]={ -16'd1108,-16'd5133,-16'd3887,16'd7448,16'd5249,-16'd4608,16'd5600,16'd2125,16'd1643,16'd2418,-16'd5891,16'd4559,-16'd3535,16'd5480,16'd1975,16'd6431,16'd4595,16'd8008,-16'd6531,16'd1418,16'd1414,16'd60,-16'd2959,16'd2102,16'd2025,-16'd3145,16'd649,16'd5757,-16'd9756,-16'd6795,16'd7310,16'd6332,-16'd6773,-16'd499,16'd2379,-16'd4478};
dout[196]={ -16'd6743,-16'd2606,16'd2513,-16'd2157,16'd7670,16'd3711,-16'd2723,16'd4070,-16'd4572,16'd3284,-16'd611,16'd893,-16'd4574,16'd3950,16'd3736,-16'd6395,16'd5590,-16'd3447,16'd1906,16'd733,16'd1575,-16'd1070,16'd3702,-16'd6364,-16'd5196,-16'd689,-16'd7165,-16'd8403,16'd4030,16'd5377,16'd7478,16'd5976,-16'd5641,-16'd6122,-16'd1297,16'd3456};
dout[197]={ 16'd5878,-16'd6944,16'd6894,-16'd3131,-16'd146,16'd4172,-16'd7148,-16'd113,-16'd6123,-16'd2040,16'd5188,16'd940,16'd275,-16'd3905,-16'd6850,-16'd5308,16'd1292,16'd1373,-16'd4674,16'd5642,-16'd6643,-16'd870,16'd5540,-16'd6,-16'd5733,16'd3096,16'd4815,16'd1282,-16'd6769,16'd6407,16'd6641,-16'd5807,16'd6601,-16'd3094,-16'd5037,-16'd4871};
dout[198]={ -16'd3114,-16'd1740,-16'd1909,16'd5594,-16'd5506,16'd3709,-16'd5335,-16'd3044,16'd1785,16'd826,-16'd878,-16'd4656,16'd118,16'd5952,16'd4408,-16'd3860,16'd4497,-16'd1031,16'd5886,-16'd3588,16'd4182,-16'd3438,-16'd1591,16'd1606,-16'd7717,16'd2562,-16'd3572,16'd3811,16'd2751,16'd7480,-16'd1167,16'd4000,16'd4775,-16'd1241,-16'd3463,-16'd5706};
dout[199]={ 16'd2536,-16'd7111,-16'd6427,-16'd4767,16'd3165,-16'd1556,-16'd3219,-16'd2573,16'd1909,-16'd503,16'd4964,16'd204,-16'd293,16'd5194,16'd645,16'd2567,-16'd4861,-16'd1224,16'd4517,-16'd4857,-16'd7885,16'd4038,16'd6158,-16'd5719,-16'd6680,16'd2386,-16'd2148,-16'd1631,16'd3892,-16'd2206,-16'd5334,16'd5054,-16'd6538,-16'd276,16'd216,-16'd2922};
dout[200]={ 16'd546,-16'd4054,-16'd1905,-16'd2215,16'd1436,16'd5131,-16'd2700,-16'd470,-16'd8014,-16'd3367,16'd5274,16'd393,16'd6135,-16'd11193,-16'd1269,16'd2609,-16'd4003,16'd11344,-16'd5152,-16'd7511,16'd3245,-16'd6492,16'd3928,16'd143,-16'd6753,16'd8302,16'd1530,-16'd6413,16'd2125,16'd734,16'd5837,-16'd3434,16'd5703,16'd2250,-16'd375,16'd3769};
dout[201]={ -16'd2329,-16'd6330,-16'd6474,-16'd6133,16'd2571,16'd4610,-16'd650,-16'd4477,-16'd1394,16'd3121,16'd7877,-16'd4550,-16'd4325,-16'd10623,-16'd3420,16'd4382,-16'd1971,-16'd1604,16'd3934,-16'd7139,-16'd6006,-16'd6691,-16'd5212,-16'd8282,-16'd9080,-16'd4294,16'd1473,-16'd5653,-16'd907,16'd612,-16'd3203,-16'd9343,-16'd5499,16'd1157,-16'd2324,-16'd6278};
dout[202]={ -16'd6833,16'd2990,16'd2471,-16'd7294,16'd3633,16'd4699,-16'd6277,16'd213,16'd2993,16'd4853,16'd3101,16'd2528,16'd2930,-16'd2765,-16'd5784,-16'd3872,-16'd7727,-16'd4801,-16'd1716,-16'd10488,16'd4428,-16'd2144,16'd6617,-16'd5808,16'd1832,16'd4112,-16'd3280,-16'd6413,16'd5853,16'd1784,16'd7830,-16'd8276,-16'd1514,16'd6950,-16'd4296,16'd3487};
dout[203]={ -16'd8705,-16'd2930,-16'd4163,16'd6214,16'd8311,-16'd4297,-16'd42,-16'd3500,16'd4091,-16'd8072,-16'd7533,-16'd1162,-16'd6649,-16'd6474,16'd7916,-16'd2902,-16'd4302,16'd6914,16'd1231,-16'd3231,16'd605,16'd1857,-16'd3874,-16'd159,-16'd7785,16'd1783,-16'd8601,16'd3192,-16'd439,16'd5935,-16'd1925,16'd6986,-16'd6835,16'd5464,-16'd14653,-16'd9184};
dout[204]={ -16'd4350,-16'd6048,-16'd1773,16'd1155,16'd4615,-16'd144,-16'd693,-16'd4179,16'd2153,16'd1819,16'd6187,16'd2870,-16'd9011,16'd3876,-16'd4807,-16'd4592,-16'd4174,16'd8768,-16'd3510,-16'd5104,-16'd1049,16'd3287,-16'd7231,-16'd4774,-16'd297,-16'd7991,-16'd2383,-16'd7718,-16'd4793,16'd851,-16'd1496,-16'd351,-16'd4316,-16'd7477,-16'd4938,-16'd248};
dout[205]={ -16'd1131,16'd8698,16'd401,-16'd3808,16'd2147,-16'd7332,-16'd2310,16'd6610,16'd4665,16'd3148,-16'd3414,-16'd4327,16'd5557,-16'd7017,16'd6033,16'd3074,16'd3967,-16'd3740,-16'd5743,-16'd3624,-16'd946,16'd2600,-16'd7255,16'd1901,-16'd10496,16'd3410,-16'd9099,-16'd5525,16'd1073,-16'd4511,16'd894,16'd3633,16'd484,16'd4805,-16'd4912,16'd5659};
dout[206]={ -16'd389,16'd4353,16'd4425,-16'd1521,-16'd2693,16'd283,-16'd3451,16'd4327,-16'd817,-16'd2713,-16'd1705,-16'd178,16'd1280,-16'd8887,16'd805,-16'd3644,16'd4805,16'd7118,16'd5636,16'd4256,16'd2891,16'd4214,16'd3655,16'd2955,-16'd3374,-16'd3787,-16'd563,16'd3372,16'd1437,16'd5944,-16'd2512,16'd4602,-16'd2961,16'd5877,-16'd10473,-16'd7021};
dout[207]={ -16'd4077,16'd579,-16'd2710,16'd4049,16'd5000,16'd2698,-16'd5840,-16'd5047,16'd2968,16'd1716,16'd3949,16'd3101,-16'd3976,16'd5988,-16'd2937,16'd2489,16'd1139,16'd3209,-16'd69,16'd2858,-16'd6932,-16'd2014,-16'd5270,-16'd5695,-16'd7954,16'd4039,16'd589,-16'd1023,16'd5467,16'd811,16'd2718,-16'd3450,-16'd5953,-16'd5918,16'd5556,16'd5876};
dout[208]={ -16'd3774,16'd1553,16'd5343,16'd1357,-16'd983,16'd7128,16'd3321,16'd451,16'd3155,-16'd6781,-16'd3690,16'd1809,16'd4465,16'd4391,16'd214,-16'd6559,16'd2760,-16'd3769,-16'd3613,16'd6739,-16'd7446,-16'd3053,16'd272,-16'd7481,-16'd8350,16'd3416,16'd6001,16'd5074,-16'd5018,16'd4635,16'd7027,16'd45,16'd1625,-16'd3692,16'd3985,16'd2841};
dout[209]={ -16'd6347,16'd624,16'd965,16'd2194,16'd1440,-16'd3439,-16'd7356,-16'd507,16'd5442,-16'd933,16'd724,-16'd6526,16'd1395,16'd4996,-16'd3656,16'd4636,-16'd4748,-16'd6447,-16'd5418,-16'd5555,-16'd5940,-16'd5926,-16'd4887,-16'd3219,-16'd5330,-16'd2734,-16'd3512,16'd2383,-16'd2786,-16'd4516,-16'd4343,-16'd8691,16'd5189,-16'd781,-16'd1827,16'd2895};
dout[210]={ -16'd2716,-16'd7602,-16'd874,16'd2248,-16'd531,16'd7803,-16'd5897,16'd1129,-16'd6840,16'd5077,16'd6139,16'd1145,-16'd491,-16'd12369,-16'd5489,-16'd6268,-16'd12155,-16'd1907,-16'd5862,-16'd7542,16'd6578,-16'd4113,16'd7448,-16'd4704,16'd1919,-16'd6342,-16'd5345,-16'd4871,16'd6298,-16'd6195,16'd2170,16'd1783,-16'd2795,16'd8247,-16'd5137,-16'd2480};
dout[211]={ -16'd6151,-16'd5593,-16'd5392,-16'd7651,16'd7840,-16'd7897,-16'd2884,-16'd4105,-16'd6033,-16'd4939,16'd1716,16'd1004,16'd4941,-16'd1957,16'd5394,16'd3779,16'd2387,16'd4851,-16'd9107,-16'd13905,-16'd304,16'd4250,16'd9239,16'd14,-16'd7390,16'd5265,16'd2939,16'd5628,16'd7803,-16'd7826,-16'd386,-16'd4319,-16'd8364,-16'd9057,16'd191,-16'd9954};
dout[212]={ -16'd4955,-16'd8840,16'd3535,16'd461,16'd3131,16'd7321,16'd2811,16'd2525,16'd1468,-16'd653,16'd3419,16'd5259,16'd4792,-16'd6881,16'd5512,16'd4193,16'd2492,16'd1367,-16'd5588,-16'd6848,16'd2645,-16'd7811,16'd3350,-16'd1852,16'd6027,16'd5250,-16'd1584,16'd2562,16'd5756,16'd4874,-16'd2589,-16'd3465,-16'd6696,16'd3834,-16'd2989,-16'd2959};
dout[213]={ 16'd3228,-16'd9535,-16'd1755,16'd3375,16'd6276,-16'd668,-16'd879,-16'd185,-16'd7800,-16'd6419,16'd1310,-16'd353,-16'd6710,-16'd2438,16'd2990,-16'd5009,-16'd7857,-16'd178,-16'd3746,-16'd3607,16'd1339,-16'd8807,-16'd3401,-16'd2115,16'd1199,-16'd94,16'd4089,16'd2891,16'd7019,16'd8876,16'd6378,-16'd5450,16'd1829,-16'd4388,-16'd5615,16'd448};
dout[214]={ -16'd1213,16'd3734,16'd3448,-16'd1195,16'd4910,-16'd6238,-16'd1160,-16'd5154,-16'd5600,-16'd6813,-16'd1822,16'd3938,-16'd2495,-16'd1766,16'd3695,16'd3347,-16'd140,16'd6060,16'd5244,16'd1727,16'd3900,16'd5227,-16'd3407,16'd638,-16'd788,-16'd6210,-16'd1738,-16'd4281,-16'd2520,16'd3176,-16'd3286,-16'd5806,-16'd6793,16'd1768,-16'd5490,16'd481};
dout[215]={ -16'd4684,16'd5868,-16'd1811,-16'd580,16'd6146,-16'd3459,16'd5878,-16'd2181,-16'd889,16'd3819,16'd2605,-16'd527,-16'd7787,-16'd2225,-16'd4527,16'd857,-16'd2449,16'd7255,16'd8223,16'd505,-16'd4298,-16'd5268,16'd4238,16'd4761,-16'd10209,16'd3334,-16'd9254,-16'd7166,-16'd5313,-16'd3368,16'd2052,16'd3142,-16'd1545,16'd5905,-16'd11233,-16'd6436};
dout[216]={ 16'd2302,-16'd7032,16'd5698,-16'd782,-16'd6003,16'd5750,16'd3305,16'd6298,16'd6624,-16'd6525,-16'd288,16'd879,16'd985,16'd5622,-16'd7263,16'd1396,16'd2285,-16'd2949,-16'd245,-16'd6657,-16'd7974,16'd2309,-16'd2158,-16'd3278,-16'd9919,16'd3915,16'd7527,-16'd4807,-16'd933,16'd4618,-16'd6203,-16'd3447,-16'd8463,-16'd5524,16'd1090,-16'd8245};
dout[217]={ 16'd3348,16'd6525,-16'd2708,-16'd3044,-16'd4703,16'd5784,16'd1490,16'd4170,-16'd4914,16'd4822,16'd5168,-16'd8523,-16'd1155,16'd2430,16'd3103,-16'd6893,16'd1025,16'd3479,16'd679,16'd27,-16'd680,16'd4040,-16'd5696,16'd6040,-16'd4801,-16'd1994,16'd7143,16'd2139,-16'd4083,16'd5176,-16'd6005,-16'd4742,-16'd4088,16'd6387,-16'd6181,16'd1822};
dout[218]={ 16'd2376,16'd7890,-16'd4689,-16'd1442,-16'd1996,-16'd5274,-16'd7607,16'd2701,-16'd3199,16'd1403,-16'd1040,16'd1426,-16'd6089,16'd2720,-16'd2243,16'd2347,16'd5944,-16'd2699,16'd6864,-16'd7854,-16'd8769,-16'd7571,16'd8285,16'd4519,-16'd8551,-16'd6477,16'd3431,-16'd6598,16'd1700,-16'd1322,-16'd1089,16'd2211,16'd3430,-16'd1641,-16'd5721,16'd3602};
dout[219]={ 16'd4748,16'd4586,16'd913,-16'd7469,-16'd6145,16'd5599,-16'd4158,-16'd3201,16'd6649,16'd4248,-16'd2879,-16'd2555,16'd3175,-16'd2746,16'd8144,16'd6656,16'd3586,-16'd5655,-16'd2273,-16'd2389,-16'd5028,-16'd4313,-16'd2269,16'd895,-16'd2856,-16'd7364,16'd3103,-16'd3864,-16'd1932,16'd3529,16'd4010,16'd330,-16'd7355,-16'd7360,16'd5635,16'd2130};
dout[220]={ -16'd177,-16'd6794,-16'd230,16'd4982,16'd7228,16'd2947,16'd848,-16'd1389,16'd3631,-16'd744,-16'd2116,16'd1138,16'd1368,-16'd6382,-16'd7961,-16'd7966,-16'd12882,16'd9852,-16'd5655,-16'd4854,-16'd3368,-16'd1049,16'd3762,16'd551,16'd3118,-16'd4585,-16'd6463,-16'd7112,16'd9902,-16'd4252,16'd2558,-16'd5116,16'd3825,16'd4341,16'd6501,-16'd9237};
dout[221]={ -16'd9357,-16'd3334,-16'd6626,-16'd8610,16'd6480,16'd1931,16'd2936,-16'd5493,16'd5381,16'd516,-16'd2218,-16'd5134,16'd6102,16'd106,16'd7209,-16'd9637,-16'd10726,16'd3424,16'd997,-16'd11147,-16'd6454,-16'd1323,16'd3998,-16'd498,-16'd2444,-16'd1489,-16'd6158,16'd2437,-16'd77,-16'd372,-16'd4170,16'd4878,-16'd6978,-16'd4223,-16'd3397,-16'd9074};
dout[222]={ -16'd4931,-16'd5109,16'd4739,-16'd6170,-16'd5841,-16'd522,-16'd6494,-16'd2295,-16'd7977,-16'd6216,16'd2502,16'd3491,16'd6742,-16'd9959,16'd8185,16'd3258,16'd1343,-16'd894,16'd1002,-16'd4803,16'd5237,16'd3207,-16'd3159,-16'd7058,-16'd4224,-16'd6881,16'd4652,-16'd4650,-16'd2375,16'd8583,16'd1778,-16'd5412,-16'd2527,-16'd5145,-16'd9201,-16'd1015};
dout[223]={ 16'd3492,16'd2033,16'd1701,-16'd7005,16'd2416,16'd1048,-16'd242,16'd820,-16'd3363,-16'd9401,16'd3906,-16'd3714,-16'd6721,16'd4028,-16'd975,-16'd5441,-16'd1704,-16'd3587,16'd5093,16'd180,-16'd1061,-16'd3205,16'd3183,-16'd229,16'd3244,16'd6066,-16'd5363,16'd2142,16'd7102,16'd5901,16'd5237,-16'd3153,-16'd5640,16'd4487,-16'd3916,16'd1659};
dout[224]={ -16'd9537,-16'd5057,-16'd4277,16'd1068,-16'd1326,16'd1809,16'd6535,-16'd6110,-16'd5179,16'd2420,-16'd1823,-16'd5438,-16'd6635,-16'd6921,-16'd3490,16'd2177,-16'd6737,-16'd2317,16'd4666,16'd4285,16'd4759,16'd1846,-16'd632,-16'd2601,16'd2395,16'd5519,-16'd7062,-16'd3012,16'd8588,16'd4764,16'd842,16'd3329,-16'd2349,16'd4601,-16'd7714,-16'd4088};
dout[225]={ -16'd572,-16'd3975,-16'd2949,16'd4191,16'd1468,16'd7398,-16'd2382,-16'd3385,16'd6228,-16'd5221,-16'd2831,-16'd8375,16'd4023,-16'd7958,-16'd2900,-16'd7244,-16'd882,16'd5662,-16'd3380,16'd169,16'd2222,16'd3543,16'd1646,-16'd4697,-16'd2837,-16'd3195,16'd3242,-16'd6987,-16'd6425,16'd4636,16'd1708,-16'd4265,-16'd3568,-16'd1802,16'd335,16'd3373};
dout[226]={ -16'd1012,16'd5183,-16'd4755,-16'd5906,-16'd101,16'd5728,-16'd5196,16'd1752,-16'd7018,-16'd3039,-16'd1616,-16'd6269,16'd4737,16'd5018,16'd1282,16'd3728,16'd6686,16'd2377,16'd2892,-16'd7468,16'd4001,-16'd1714,-16'd4133,16'd4310,16'd5678,-16'd2255,16'd3091,-16'd5800,-16'd2658,-16'd1450,16'd3906,16'd4105,16'd348,16'd3457,-16'd10178,-16'd808};
dout[227]={ 16'd4760,16'd7526,-16'd5369,-16'd4776,16'd444,16'd5948,-16'd1016,16'd3815,16'd6720,-16'd2385,-16'd544,-16'd6908,-16'd451,-16'd1553,-16'd1075,16'd6871,16'd3197,-16'd3021,16'd2193,16'd955,16'd7119,-16'd127,16'd2227,-16'd1156,16'd3363,16'd708,-16'd116,16'd5155,-16'd3162,-16'd5369,-16'd2845,-16'd9222,16'd1662,-16'd1812,-16'd8443,-16'd5975};
dout[228]={ -16'd4551,-16'd850,16'd3627,16'd334,16'd6012,16'd890,-16'd2649,-16'd2204,16'd3429,-16'd8889,16'd4047,-16'd8026,-16'd1447,16'd4454,-16'd2841,16'd6182,16'd949,-16'd2341,16'd5047,-16'd1172,-16'd5059,-16'd3546,16'd2236,16'd5913,-16'd8720,16'd251,16'd5395,-16'd3418,-16'd37,-16'd4502,-16'd3368,16'd3260,-16'd2246,16'd6686,16'd3302,-16'd5807};
dout[229]={ 16'd6,16'd4644,16'd2993,-16'd3819,-16'd3388,-16'd607,16'd2653,-16'd3661,16'd1969,-16'd884,16'd1336,16'd2804,-16'd2964,-16'd4264,-16'd2207,16'd452,16'd3014,-16'd8526,16'd5409,-16'd7909,-16'd101,-16'd4760,-16'd6971,-16'd445,-16'd4225,16'd1662,-16'd8659,16'd5553,16'd5073,16'd2869,16'd1711,-16'd6793,16'd5703,-16'd2093,16'd4554,-16'd936};
dout[230]={ 16'd7638,-16'd3885,-16'd1925,-16'd5625,16'd6483,-16'd237,-16'd3147,-16'd708,-16'd706,-16'd6322,-16'd1022,-16'd1548,16'd1097,-16'd2080,-16'd5228,-16'd2458,-16'd667,16'd4258,-16'd2914,-16'd6212,16'd5606,-16'd2034,-16'd576,16'd6260,16'd3646,16'd3135,-16'd9208,16'd1792,16'd4708,16'd2725,-16'd6725,-16'd4029,-16'd5497,16'd12357,-16'd4904,-16'd874};
dout[231]={ 16'd730,16'd4948,16'd1351,-16'd5879,-16'd338,-16'd3341,-16'd415,-16'd1127,16'd3068,16'd1450,16'd1220,16'd1693,16'd5477,-16'd10308,16'd523,-16'd8245,-16'd9869,-16'd6528,-16'd7601,-16'd7143,16'd6180,-16'd2994,-16'd3092,-16'd8636,16'd2788,-16'd5610,16'd1395,-16'd1876,-16'd1666,-16'd2384,-16'd554,16'd368,-16'd675,16'd2409,-16'd3817,-16'd3440};
dout[232]={ -16'd9549,-16'd6793,-16'd4621,-16'd2271,16'd330,16'd2134,16'd1999,-16'd9257,-16'd7159,16'd2724,-16'd832,-16'd2634,16'd630,16'd2396,16'd7015,-16'd2736,-16'd7259,-16'd3186,16'd4083,-16'd7675,16'd1607,16'd8953,16'd2648,-16'd9391,-16'd5813,-16'd1638,16'd1492,16'd6307,16'd222,16'd3767,-16'd1946,-16'd9272,-16'd3521,-16'd4317,-16'd7123,16'd528};
dout[233]={ -16'd4200,16'd5031,-16'd5530,16'd2336,16'd1169,-16'd10,-16'd7729,-16'd6347,16'd1644,16'd1764,16'd4139,-16'd1555,16'd1086,16'd1859,16'd6266,-16'd5955,-16'd7237,-16'd8080,16'd4987,-16'd1684,-16'd2744,-16'd5124,16'd4364,16'd3379,16'd2211,-16'd6372,-16'd7545,16'd3190,-16'd3829,16'd9500,-16'd2039,16'd1800,-16'd6598,-16'd1764,16'd2055,-16'd3828};
dout[234]={ -16'd7672,-16'd5101,16'd1753,16'd5758,16'd6029,16'd1539,16'd7085,16'd472,-16'd5413,-16'd3535,-16'd7596,-16'd6613,-16'd4244,16'd530,-16'd7612,-16'd3703,16'd4806,-16'd15,-16'd4367,-16'd786,-16'd3723,-16'd993,16'd8546,-16'd3851,-16'd1224,-16'd3142,-16'd6734,16'd2776,-16'd1500,-16'd873,-16'd6630,-16'd244,-16'd1430,16'd612,-16'd458,16'd5308};
dout[235]={ 16'd6409,-16'd2202,-16'd6392,16'd704,16'd5244,16'd3033,-16'd4636,16'd3752,-16'd3209,-16'd1424,-16'd2833,16'd4170,16'd3902,16'd2803,-16'd7795,-16'd621,16'd7033,16'd1210,16'd8564,-16'd4006,16'd5322,-16'd137,-16'd4792,16'd4093,-16'd4192,16'd1873,-16'd5496,16'd6912,16'd3469,16'd3031,16'd5176,16'd421,16'd1245,-16'd3653,-16'd7662,16'd3531};
dout[236]={ -16'd6573,16'd3855,-16'd2185,-16'd1459,-16'd3140,16'd896,16'd5877,-16'd5590,-16'd5489,-16'd2661,16'd2928,-16'd3438,-16'd3527,-16'd3940,16'd3680,-16'd181,-16'd7,16'd6802,-16'd132,16'd6047,16'd5020,16'd6532,16'd6735,16'd4918,-16'd2923,16'd5844,-16'd3924,16'd104,16'd2476,16'd6985,16'd2919,-16'd1458,16'd3708,-16'd1359,-16'd10898,16'd3781};
dout[237]={ 16'd5470,-16'd6946,-16'd7038,-16'd3444,-16'd2962,-16'd1417,16'd3301,16'd4687,16'd5850,-16'd1107,-16'd2187,-16'd3232,16'd1523,16'd3919,-16'd2105,-16'd1983,-16'd2744,16'd1694,-16'd1821,16'd3530,-16'd1256,16'd2516,-16'd6448,-16'd5438,-16'd5035,16'd4551,16'd6932,16'd5698,16'd3022,-16'd5236,-16'd5084,-16'd5871,16'd6471,16'd1479,-16'd7625,16'd3940};
dout[238]={ 16'd4636,16'd847,-16'd3864,16'd3210,16'd6027,-16'd5321,-16'd4601,16'd1362,16'd404,-16'd764,16'd4812,-16'd7834,16'd166,16'd3252,16'd534,-16'd5554,-16'd1313,-16'd3565,16'd317,-16'd8846,-16'd364,16'd4319,16'd7265,16'd6386,16'd3601,-16'd5889,-16'd3943,-16'd3221,-16'd987,16'd5904,16'd5945,16'd4105,-16'd3670,16'd1783,16'd3399,-16'd4405};
dout[239]={ 16'd4198,-16'd3072,16'd765,-16'd3707,-16'd245,-16'd5064,16'd4291,16'd1372,16'd5423,16'd1539,16'd2030,16'd5006,16'd4345,16'd600,-16'd286,16'd3010,-16'd1383,-16'd920,16'd6259,-16'd8011,-16'd8033,16'd2072,-16'd4013,16'd1062,-16'd4570,-16'd3528,-16'd7202,16'd549,-16'd2091,16'd2515,16'd1981,-16'd1089,-16'd5397,-16'd5908,-16'd9320,-16'd2037};
dout[240]={ -16'd1058,16'd4774,16'd3484,-16'd4546,-16'd4338,16'd6451,16'd1877,16'd763,16'd4368,-16'd5050,16'd3210,-16'd5987,-16'd4439,-16'd11973,16'd1508,-16'd2519,-16'd88,16'd1208,-16'd11533,16'd1110,16'd586,16'd5277,-16'd267,16'd2176,16'd3692,-16'd3957,-16'd4250,16'd4912,16'd991,16'd3504,16'd2593,-16'd5222,-16'd1287,16'd11168,-16'd1158,-16'd12675};
dout[241]={ -16'd6471,-16'd7382,-16'd6078,16'd6605,-16'd6240,-16'd7232,-16'd7499,-16'd4009,-16'd1524,16'd3476,-16'd886,16'd3133,16'd1651,-16'd5065,-16'd4846,16'd2411,-16'd1093,16'd239,-16'd1823,-16'd3229,-16'd4835,16'd7123,16'd66,-16'd224,-16'd9695,16'd1143,-16'd3442,16'd4120,-16'd2458,16'd4411,16'd2408,-16'd212,16'd5699,16'd1937,-16'd4678,-16'd1497};
dout[242]={ -16'd138,-16'd1010,16'd4192,-16'd3955,-16'd4648,-16'd2078,-16'd2763,16'd2865,-16'd5117,-16'd3834,-16'd1271,-16'd40,16'd5478,-16'd4345,-16'd6478,-16'd4383,-16'd6481,16'd1496,-16'd8080,-16'd5111,16'd4166,16'd8799,16'd5649,16'd1659,16'd5315,-16'd7978,16'd3464,16'd2806,16'd10155,16'd3192,-16'd7215,-16'd2345,16'd4669,16'd5410,-16'd1433,-16'd8718};
dout[243]={ -16'd7754,-16'd6206,-16'd3861,16'd6567,-16'd2919,-16'd2469,-16'd2653,-16'd4040,-16'd2287,-16'd10128,16'd1719,-16'd2344,16'd5986,16'd4802,-16'd4776,16'd2497,-16'd4999,-16'd1051,-16'd5696,-16'd4559,16'd7313,16'd1084,-16'd571,16'd4806,16'd6433,-16'd229,16'd1058,-16'd64,16'd8986,16'd1894,-16'd3893,16'd4838,-16'd1159,16'd4765,-16'd9252,-16'd2268};
dout[244]={ 16'd5095,-16'd7325,16'd6003,-16'd3238,-16'd5692,16'd6032,-16'd2094,-16'd8208,-16'd5835,-16'd343,16'd5311,-16'd1765,16'd4348,-16'd2318,-16'd323,-16'd5681,16'd3982,-16'd1685,16'd7245,-16'd1542,-16'd925,-16'd3662,16'd5334,16'd4758,16'd3926,-16'd6285,-16'd5111,-16'd6456,-16'd2623,16'd5585,16'd1007,-16'd2427,16'd802,-16'd7143,-16'd6025,-16'd2426};
dout[245]={ 16'd2023,16'd3301,-16'd1126,-16'd1880,-16'd2962,-16'd6993,-16'd3523,16'd7123,-16'd3642,-16'd8254,-16'd5022,-16'd6160,16'd6920,16'd5026,-16'd655,16'd2386,-16'd1501,-16'd2045,-16'd1439,16'd6481,16'd1895,16'd5096,-16'd1680,-16'd6061,-16'd6241,-16'd1465,-16'd3575,-16'd1862,-16'd4777,-16'd5582,-16'd6828,-16'd425,16'd4706,-16'd3821,-16'd9610,16'd1301};
dout[246]={ 16'd1998,16'd2066,16'd3371,16'd6886,-16'd7341,16'd3990,-16'd717,16'd1321,-16'd4100,-16'd4172,-16'd1116,-16'd5751,-16'd2084,16'd367,-16'd7216,-16'd6874,16'd2987,16'd488,16'd4906,-16'd4772,-16'd1884,16'd1905,16'd5226,16'd3038,-16'd2106,-16'd5730,-16'd6991,16'd5087,-16'd7302,16'd433,16'd1018,-16'd6109,-16'd4773,-16'd7156,16'd2282,-16'd4316};
dout[247]={ 16'd944,-16'd7888,16'd7310,-16'd3574,-16'd4663,16'd1059,-16'd3787,-16'd4239,-16'd1012,-16'd2983,-16'd2921,-16'd2299,-16'd5657,16'd3492,16'd3781,16'd1268,-16'd672,-16'd2532,-16'd5195,-16'd2984,-16'd1312,-16'd2457,16'd2458,-16'd3853,-16'd3541,16'd2721,16'd4625,-16'd8011,16'd5574,-16'd2330,-16'd5492,16'd862,-16'd4808,-16'd4721,-16'd8125,16'd357};
dout[248]={ 16'd5649,16'd2957,16'd497,16'd982,16'd7241,16'd1785,16'd282,-16'd1428,-16'd136,-16'd4913,-16'd8330,-16'd427,-16'd4602,-16'd5568,-16'd1429,16'd4249,16'd4015,-16'd6390,-16'd7391,16'd8092,-16'd2649,16'd3951,-16'd7041,-16'd409,-16'd5583,16'd3344,-16'd22,16'd2802,-16'd4731,16'd3181,16'd5063,16'd2610,-16'd5054,-16'd5268,16'd759,-16'd1775};
dout[249]={ -16'd814,16'd3321,16'd2440,-16'd1647,16'd4359,-16'd138,-16'd1414,-16'd2531,-16'd5871,16'd4374,-16'd3178,16'd1994,16'd5187,-16'd4194,16'd1768,-16'd32,-16'd5702,-16'd5740,-16'd951,16'd5836,16'd6967,16'd3658,16'd1277,16'd9059,16'd4451,-16'd663,16'd2020,16'd6580,-16'd3852,-16'd6532,16'd2762,-16'd4065,16'd3384,-16'd8770,-16'd4654,16'd2714};
dout[250]={ 16'd8990,16'd4728,-16'd9335,16'd3811,-16'd10625,-16'd4699,-16'd4983,-16'd8348,-16'd7100,-16'd768,16'd2864,16'd2726,-16'd1265,-16'd3398,-16'd1495,-16'd5904,16'd3584,-16'd2540,-16'd281,-16'd1101,-16'd4171,16'd8351,-16'd199,-16'd2281,16'd2684,16'd5561,-16'd6670,16'd1325,16'd1825,-16'd4850,-16'd5971,-16'd2560,16'd9772,16'd14038,16'd3167,-16'd1100};
dout[251]={ -16'd2806,16'd1628,16'd2312,16'd533,16'd2174,16'd1719,-16'd995,-16'd3501,-16'd5219,16'd2771,-16'd3705,-16'd7708,16'd4313,-16'd8022,16'd5667,-16'd3380,-16'd394,-16'd5360,-16'd1566,-16'd933,-16'd4310,-16'd795,-16'd3391,16'd883,16'd584,-16'd3499,16'd2599,-16'd3693,-16'd2639,16'd4927,16'd5614,-16'd1958,16'd7174,-16'd6612,16'd2607,-16'd11362};
dout[252]={ -16'd1910,-16'd6453,16'd92,-16'd3723,-16'd12672,-16'd4228,16'd6383,-16'd5853,16'd737,-16'd8481,-16'd2079,-16'd3635,16'd2509,16'd575,16'd1735,-16'd777,-16'd1677,-16'd4516,-16'd1586,-16'd4383,-16'd1782,16'd535,16'd2746,-16'd3937,-16'd2422,16'd3284,-16'd2971,-16'd7620,16'd7488,16'd3053,-16'd7330,-16'd1638,-16'd6157,16'd1119,-16'd768,-16'd6377};
dout[253]={ -16'd4178,16'd1492,-16'd3685,-16'd5539,-16'd3487,-16'd62,-16'd3571,-16'd27,-16'd3885,-16'd5025,16'd3098,-16'd1363,-16'd2222,16'd1536,-16'd9966,-16'd7975,16'd4684,-16'd15,16'd1924,-16'd1764,16'd1045,16'd10033,16'd7232,-16'd897,-16'd920,16'd4785,-16'd6728,-16'd724,16'd7133,16'd8008,16'd2364,-16'd5518,-16'd3246,-16'd274,-16'd8952,16'd2172};
dout[254]={ -16'd514,-16'd3908,-16'd3824,16'd3322,-16'd6711,-16'd2994,16'd7189,-16'd6915,-16'd8182,-16'd719,16'd2107,16'd5537,-16'd2479,-16'd394,-16'd4654,16'd5858,16'd7528,16'd1651,-16'd4449,-16'd5140,16'd2097,-16'd2389,-16'd5700,-16'd1505,-16'd5186,-16'd2543,16'd3403,-16'd3104,16'd1632,-16'd582,16'd4226,-16'd4303,16'd6970,-16'd2885,16'd4165,16'd5382};
dout[255]={ 16'd1281,16'd3959,-16'd7069,16'd6124,-16'd5789,-16'd7429,-16'd4318,16'd453,-16'd6344,16'd177,-16'd2541,-16'd4109,-16'd5974,-16'd1860,-16'd771,-16'd7057,-16'd2600,16'd1031,-16'd2196,-16'd443,16'd3490,16'd2475,16'd1943,-16'd5489,16'd3459,-16'd6449,-16'd1551,-16'd6557,-16'd7089,16'd5066,-16'd1354,-16'd211,-16'd6393,-16'd6079,16'd3578,-16'd245};
dout[256]={ 16'd5670,16'd1635,-16'd3586,-16'd3590,16'd6312,-16'd5612,-16'd6168,16'd1115,-16'd3152,-16'd6550,-16'd5352,-16'd3751,16'd2078,16'd5145,16'd7320,16'd2329,16'd4421,16'd866,16'd190,16'd7339,16'd662,16'd2956,-16'd5567,-16'd4730,-16'd6913,-16'd7562,16'd1307,16'd3364,-16'd4169,-16'd6491,-16'd4920,16'd1949,16'd5270,-16'd2500,16'd5031,-16'd573};
dout[257]={ 16'd3372,16'd3637,16'd2822,-16'd2070,-16'd4994,-16'd4935,-16'd4106,16'd3684,-16'd5702,16'd1427,-16'd3275,16'd3978,16'd5785,16'd1969,16'd7797,-16'd2704,16'd6642,-16'd3553,16'd2024,16'd6734,16'd2754,16'd200,-16'd3789,-16'd5467,-16'd6847,-16'd7556,-16'd727,-16'd985,-16'd1122,16'd7645,-16'd4055,-16'd591,16'd4060,16'd4960,-16'd4962,-16'd633};
dout[258]={ 16'd641,-16'd5403,16'd1524,16'd2614,16'd3830,16'd1586,-16'd7164,16'd944,-16'd7398,-16'd5445,-16'd4387,-16'd7306,16'd2338,-16'd6545,-16'd3237,16'd3236,16'd2935,16'd5550,16'd2031,16'd5567,-16'd7879,16'd2866,-16'd4095,16'd5893,16'd8000,-16'd6228,-16'd5130,-16'd7978,-16'd5467,16'd4435,-16'd7387,-16'd3313,-16'd3921,16'd4660,-16'd2167,16'd4258};
dout[259]={ 16'd781,-16'd8532,16'd80,-16'd4935,16'd4025,16'd3567,16'd509,16'd7732,-16'd2673,16'd3641,16'd1283,-16'd6722,16'd5817,16'd3301,-16'd4179,-16'd8010,-16'd5228,16'd6001,16'd435,16'd6529,-16'd2511,16'd6089,-16'd5373,16'd4322,-16'd5528,16'd3501,-16'd4268,-16'd948,16'd6239,16'd1190,-16'd2239,-16'd726,-16'd6012,-16'd4476,-16'd5446,16'd6742};
dout[260]={ -16'd4888,-16'd1627,-16'd5882,-16'd3751,-16'd7575,16'd6449,16'd2009,-16'd1720,-16'd3132,16'd2815,-16'd5287,16'd3229,-16'd1556,-16'd6609,16'd3368,-16'd4086,-16'd2870,16'd6228,-16'd8,16'd3266,16'd6046,-16'd4958,-16'd4266,-16'd3126,16'd3603,16'd5762,16'd2591,-16'd5063,16'd5833,16'd5233,-16'd943,16'd3032,-16'd1375,16'd5096,16'd3838,-16'd12079};
dout[261]={ 16'd2640,16'd3298,16'd2503,16'd7927,-16'd393,16'd4474,-16'd4293,-16'd2042,16'd5942,-16'd7269,16'd1605,16'd4506,-16'd3023,-16'd6853,16'd2824,16'd1943,-16'd7718,16'd2451,-16'd4299,-16'd3257,16'd6828,16'd777,-16'd4365,-16'd9291,-16'd7041,-16'd7577,-16'd4188,16'd2362,-16'd4611,16'd5345,16'd4475,16'd4864,-16'd247,-16'd5031,-16'd3901,-16'd324};
dout[262]={ -16'd7,-16'd7511,-16'd1812,16'd4697,-16'd3605,16'd4772,16'd3883,-16'd335,-16'd2035,-16'd3308,16'd4408,16'd595,-16'd697,-16'd425,16'd4450,16'd3737,-16'd5584,16'd6683,-16'd4333,16'd5425,-16'd7303,16'd2418,16'd5118,16'd188,16'd4643,-16'd310,16'd691,16'd4963,16'd5538,-16'd2613,-16'd1371,16'd4848,-16'd43,-16'd3265,-16'd4396,-16'd5872};
dout[263]={ 16'd6248,-16'd1900,16'd8308,-16'd4293,-16'd3726,-16'd1032,-16'd3014,-16'd1306,-16'd3756,16'd3924,-16'd7640,-16'd2355,16'd768,16'd137,-16'd3014,16'd4077,-16'd5385,-16'd557,16'd6449,-16'd1921,-16'd5154,-16'd4808,-16'd3199,-16'd2062,16'd5791,-16'd6889,16'd4323,16'd5588,16'd4385,-16'd2945,16'd2659,16'd4169,-16'd4657,16'd4959,-16'd732,-16'd491};
dout[264]={ -16'd4067,16'd4296,16'd6098,16'd6932,-16'd3194,16'd6141,-16'd6558,-16'd6766,-16'd7684,-16'd8589,16'd2100,16'd2355,16'd2852,-16'd6923,-16'd7782,-16'd5374,16'd3157,-16'd6129,-16'd2611,16'd5909,16'd809,16'd4974,16'd273,-16'd3412,-16'd1988,16'd2558,-16'd7360,-16'd8437,16'd2542,16'd492,16'd5341,-16'd1566,16'd2736,-16'd6939,-16'd3171,16'd2934};
dout[265]={ 16'd215,-16'd6139,16'd6357,-16'd1340,16'd2992,-16'd3053,16'd5401,16'd175,16'd4552,-16'd3734,16'd1484,-16'd4302,16'd3888,-16'd5167,-16'd5523,16'd1625,-16'd1244,16'd12,-16'd7062,16'd1341,-16'd8475,16'd327,-16'd6198,-16'd8752,16'd220,16'd5906,16'd2139,-16'd6520,16'd894,-16'd7287,-16'd5186,-16'd7126,16'd763,-16'd1091,-16'd5228,-16'd2234};
dout[266]={ 16'd2757,-16'd856,-16'd651,-16'd4269,-16'd3431,16'd2890,16'd2665,-16'd475,-16'd4814,16'd2095,16'd5548,16'd5258,16'd274,16'd6503,16'd1999,-16'd2032,-16'd5617,-16'd4926,16'd5434,-16'd1559,16'd5170,-16'd6112,16'd6114,-16'd1393,16'd1125,16'd5381,-16'd8087,-16'd367,-16'd1251,16'd1412,-16'd5918,16'd3980,16'd3189,16'd6044,-16'd4977,16'd3738};
dout[267]={ -16'd5624,-16'd6206,-16'd6809,16'd5196,16'd3984,-16'd1754,-16'd3236,16'd4187,16'd4191,16'd4922,-16'd878,16'd2995,-16'd6484,-16'd4461,16'd1697,-16'd1036,-16'd4303,-16'd819,-16'd4858,16'd6733,16'd4974,16'd5156,16'd939,16'd1675,-16'd5948,16'd6746,-16'd1202,16'd2046,-16'd5442,16'd4078,-16'd5497,16'd5482,16'd139,16'd6430,16'd2426,16'd677};
dout[268]={ 16'd5973,16'd2771,16'd2582,16'd4964,-16'd421,16'd5855,-16'd3945,-16'd664,16'd5694,-16'd5556,-16'd173,16'd3888,16'd415,16'd1113,-16'd1779,16'd7651,-16'd4276,16'd3951,-16'd6942,16'd6351,16'd4265,-16'd7776,16'd5795,16'd3911,-16'd720,-16'd2970,-16'd5699,-16'd479,-16'd6863,-16'd4363,-16'd6719,-16'd5350,16'd5566,16'd902,16'd3350,-16'd2954};
dout[269]={ 16'd4061,-16'd4931,-16'd4029,16'd2008,-16'd425,-16'd3812,16'd1807,16'd6171,-16'd174,-16'd1838,-16'd808,-16'd3385,-16'd2525,-16'd7267,16'd4758,-16'd1333,-16'd4268,-16'd75,16'd680,16'd4975,-16'd1825,16'd5357,-16'd3414,-16'd3539,-16'd960,16'd4392,16'd851,-16'd7355,-16'd107,-16'd1570,-16'd2898,16'd1359,-16'd5081,16'd3900,-16'd7238,16'd3181};
dout[270]={ 16'd4477,16'd3389,-16'd6629,16'd2393,16'd3101,-16'd3572,-16'd2269,16'd4109,-16'd1180,-16'd750,16'd3999,16'd2903,-16'd2881,-16'd5285,16'd6390,16'd2257,16'd1812,16'd2238,-16'd3790,-16'd7543,16'd5246,16'd1360,16'd1363,16'd6461,16'd1123,-16'd3155,16'd2818,16'd1006,16'd10246,16'd1393,-16'd6785,-16'd2878,-16'd371,16'd7708,-16'd9022,-16'd7246};
dout[271]={ -16'd2231,16'd4680,-16'd7122,16'd5321,-16'd748,-16'd7832,-16'd5817,16'd3870,16'd5553,16'd2469,16'd4512,16'd1593,-16'd12589,-16'd563,-16'd1429,-16'd6245,16'd131,16'd8227,-16'd1107,-16'd438,-16'd2254,16'd5841,-16'd3368,-16'd4693,16'd553,16'd167,-16'd8691,-16'd5808,16'd1386,16'd1162,-16'd29,16'd476,16'd7165,16'd7967,16'd2795,16'd1263};
dout[272]={ 16'd3294,-16'd428,-16'd180,-16'd7211,-16'd2348,16'd1576,16'd73,-16'd9985,-16'd1329,-16'd3176,16'd2217,16'd4487,16'd2135,-16'd8769,-16'd6102,-16'd532,16'd2909,16'd2942,16'd5808,16'd1490,16'd7711,-16'd7030,-16'd7002,-16'd4085,-16'd3902,16'd1709,-16'd9689,-16'd306,-16'd210,-16'd6132,16'd2150,-16'd3199,-16'd6692,-16'd8655,-16'd2375,-16'd8228};
dout[273]={ 16'd6268,-16'd4534,16'd7429,16'd6424,16'd2360,-16'd3756,16'd3264,-16'd5048,16'd6136,16'd31,-16'd8934,16'd619,-16'd1489,-16'd3697,-16'd7271,-16'd5027,-16'd2795,-16'd4388,16'd1596,-16'd4520,16'd4431,16'd4049,16'd2808,-16'd1882,-16'd4675,-16'd3307,16'd3105,-16'd6816,-16'd2096,-16'd7675,16'd5938,-16'd1603,16'd3648,16'd6519,-16'd6252,-16'd4710};
dout[274]={ -16'd311,-16'd1181,16'd1912,16'd435,-16'd3662,16'd4651,-16'd3518,-16'd973,-16'd518,16'd55,16'd5061,16'd5206,-16'd5437,-16'd6094,-16'd6099,-16'd1939,16'd765,-16'd6961,16'd5138,-16'd6794,-16'd532,16'd5233,16'd2003,16'd2708,-16'd3942,-16'd1012,16'd5941,-16'd5315,16'd1712,16'd4886,16'd2782,-16'd7684,16'd1638,-16'd877,-16'd3868,-16'd1357};
dout[275]={ -16'd3232,16'd5405,16'd5558,16'd5821,16'd4061,-16'd4576,-16'd2196,16'd635,-16'd3384,-16'd205,16'd5802,-16'd7131,16'd5863,-16'd2880,-16'd5472,-16'd6350,-16'd4998,-16'd5744,16'd4116,16'd6026,16'd4273,16'd6049,16'd7274,16'd4877,16'd3804,-16'd230,-16'd3583,-16'd5300,16'd4169,-16'd2817,-16'd2402,-16'd7784,-16'd5465,-16'd2761,16'd4033,-16'd4038};
dout[276]={ 16'd2285,-16'd8308,16'd3432,16'd3164,16'd2037,16'd2079,-16'd2908,16'd1259,-16'd4482,-16'd436,-16'd6433,16'd4742,-16'd5723,-16'd1261,-16'd5249,16'd4156,16'd498,-16'd2414,16'd2266,-16'd6002,16'd6469,16'd6524,16'd533,16'd580,16'd6438,-16'd800,-16'd1651,16'd5380,-16'd5396,-16'd5706,16'd1169,16'd4487,-16'd284,-16'd2646,16'd4695,16'd1214};
dout[277]={ 16'd2521,-16'd844,16'd1229,16'd1805,16'd6409,-16'd472,-16'd5639,16'd2192,16'd5514,16'd1494,-16'd1356,-16'd6186,-16'd3525,-16'd3361,-16'd4538,16'd7046,16'd1302,16'd4704,-16'd5949,-16'd6073,-16'd1416,-16'd1152,-16'd6843,16'd4351,-16'd745,16'd6301,-16'd5166,16'd2847,16'd2634,-16'd6482,16'd3040,-16'd2154,-16'd1003,-16'd6720,-16'd7454,-16'd958};
dout[278]={ -16'd643,-16'd5595,16'd4986,-16'd5028,-16'd1289,-16'd6727,16'd2843,16'd5961,16'd1090,-16'd4992,16'd6944,-16'd294,-16'd3853,16'd2213,-16'd1828,-16'd4373,16'd7588,16'd3629,-16'd1071,-16'd2734,16'd6853,-16'd6901,16'd5221,16'd3776,-16'd639,-16'd5214,16'd2333,-16'd6618,-16'd6541,-16'd5693,16'd7104,16'd3799,-16'd1418,-16'd8077,-16'd6947,16'd3016};
dout[279]={ -16'd7040,16'd6568,-16'd4253,-16'd2237,-16'd6839,16'd7359,16'd1931,16'd1096,16'd7904,-16'd1184,16'd5854,16'd1697,16'd2794,-16'd4970,16'd6526,16'd1609,16'd2128,16'd6957,16'd2207,-16'd5716,-16'd2658,-16'd208,16'd6693,-16'd329,-16'd731,-16'd4554,-16'd792,-16'd2877,-16'd4984,16'd4574,16'd1423,16'd3582,-16'd2737,16'd3519,16'd5770,16'd7382};
dout[280]={ 16'd7877,16'd4260,-16'd4593,16'd302,-16'd9441,-16'd1427,16'd6656,-16'd7909,-16'd1256,-16'd4951,-16'd6697,-16'd857,-16'd8192,16'd1807,-16'd2972,16'd7656,-16'd2378,16'd3555,16'd5737,-16'd7586,-16'd429,16'd3961,-16'd7314,-16'd2368,16'd5409,16'd8706,-16'd2876,-16'd4491,16'd3889,-16'd2682,-16'd144,16'd3189,16'd1384,16'd10019,16'd5059,-16'd349};
dout[281]={ -16'd3086,16'd2347,16'd1010,-16'd2214,-16'd10076,16'd4078,16'd1186,-16'd6445,16'd4145,-16'd1244,-16'd1488,-16'd5283,-16'd1602,-16'd5113,-16'd5517,16'd4252,-16'd4357,16'd3153,16'd6296,-16'd1015,16'd3757,-16'd3794,16'd2365,-16'd3239,-16'd1541,-16'd1209,16'd61,-16'd5956,16'd3359,16'd2593,-16'd3200,16'd2781,16'd2472,16'd236,-16'd6407,16'd750};
dout[282]={ -16'd6401,16'd5373,-16'd4275,16'd6436,16'd472,-16'd259,-16'd4134,-16'd8269,16'd1594,16'd7204,-16'd6079,-16'd872,16'd2220,16'd5214,16'd3397,-16'd6949,-16'd3192,-16'd3426,-16'd2372,16'd644,-16'd3901,-16'd2483,16'd6241,16'd1772,16'd2235,-16'd4878,-16'd455,-16'd3441,-16'd4735,-16'd776,16'd4698,-16'd3752,-16'd1016,-16'd4450,16'd4103,-16'd2552};
dout[283]={ 16'd2673,16'd1940,-16'd7340,16'd4637,16'd592,-16'd7334,16'd7912,16'd3558,-16'd1066,16'd4275,-16'd8125,16'd4582,-16'd2507,-16'd3976,-16'd7707,16'd888,-16'd1151,16'd2839,16'd9469,16'd1075,-16'd1141,16'd336,16'd5828,-16'd6649,16'd3892,16'd387,16'd4267,16'd591,-16'd4714,-16'd7340,16'd5474,-16'd6829,-16'd6323,16'd397,16'd5674,16'd6179};
dout[284]={ -16'd4725,16'd5436,-16'd3585,16'd3665,-16'd1210,16'd1242,16'd3766,-16'd2228,-16'd7939,16'd6634,16'd2339,16'd3362,-16'd568,16'd3249,16'd8944,16'd1771,16'd3062,-16'd2340,-16'd798,16'd6390,-16'd4518,16'd4175,16'd6296,-16'd8375,16'd2248,16'd4081,-16'd7660,-16'd1339,16'd5575,16'd6938,16'd5813,16'd876,16'd4685,16'd193,16'd116,-16'd620};
dout[285]={ -16'd4414,-16'd2144,16'd2187,16'd1863,16'd5298,16'd4731,-16'd6879,-16'd1722,-16'd7984,16'd1122,16'd3937,-16'd1065,-16'd2129,-16'd1144,16'd5280,-16'd696,16'd5036,-16'd6471,16'd5842,16'd5275,16'd3331,16'd1601,-16'd135,16'd5424,-16'd545,-16'd4179,16'd6793,-16'd7886,16'd1173,-16'd1461,-16'd1642,16'd2237,-16'd2301,-16'd264,-16'd449,16'd5888};
dout[286]={ -16'd790,-16'd698,16'd7080,-16'd1777,16'd1936,-16'd3973,-16'd5558,16'd477,16'd3111,16'd3023,-16'd5595,16'd6316,16'd6651,-16'd7564,16'd696,-16'd2433,16'd2175,16'd4966,-16'd1080,16'd2026,-16'd7060,-16'd7107,-16'd4888,-16'd2785,-16'd5449,-16'd3498,16'd4842,-16'd7056,-16'd5319,-16'd8173,-16'd4347,16'd4695,-16'd5245,16'd6263,-16'd7494,-16'd5238};
dout[287]={ 16'd86,-16'd687,16'd1008,16'd6683,16'd1647,-16'd5506,16'd1160,16'd7421,-16'd2509,-16'd54,16'd1059,-16'd5202,-16'd995,16'd4479,16'd1866,16'd3939,-16'd6404,16'd5164,-16'd4717,-16'd4806,-16'd6761,16'd3010,-16'd519,16'd3673,-16'd4305,-16'd3816,16'd6041,16'd3340,16'd2647,16'd423,-16'd3422,16'd2825,16'd3244,-16'd7337,16'd2992,-16'd2908};
dout[288]={ -16'd1225,-16'd1010,-16'd317,16'd2921,-16'd6150,-16'd204,-16'd9277,-16'd4011,16'd5629,16'd552,-16'd3478,-16'd3187,-16'd2242,16'd3342,16'd4869,-16'd905,16'd3539,16'd5510,-16'd6545,-16'd1399,-16'd3256,-16'd4223,16'd2163,16'd487,-16'd4428,-16'd32,16'd5422,16'd691,-16'd6252,16'd4395,-16'd2597,16'd6679,16'd1200,-16'd8407,-16'd7655,16'd5157};
dout[289]={ 16'd2981,-16'd3579,-16'd3098,16'd6551,16'd6761,16'd5820,16'd1923,-16'd3355,16'd2288,16'd4908,16'd7450,16'd5424,-16'd5184,16'd4257,16'd1291,16'd3764,16'd2904,-16'd3806,16'd6359,16'd1992,16'd2781,-16'd7064,-16'd3782,-16'd280,16'd4688,16'd618,16'd428,16'd314,16'd1571,16'd5702,16'd17,-16'd6649,-16'd431,-16'd5665,-16'd104,16'd4291};
dout[290]={ -16'd1312,16'd3082,16'd2240,-16'd8589,16'd543,-16'd1929,-16'd146,16'd4372,-16'd2903,16'd2530,-16'd1892,-16'd2953,-16'd10665,-16'd10619,-16'd4435,-16'd6791,-16'd7571,16'd8561,-16'd2167,-16'd3408,16'd10114,-16'd6771,16'd3306,-16'd6087,-16'd5616,-16'd6328,-16'd11086,16'd964,16'd4172,-16'd3060,-16'd1351,16'd7750,16'd1187,16'd2725,-16'd1636,-16'd2538};
dout[291]={ -16'd708,-16'd5881,16'd2006,-16'd2101,-16'd5602,16'd3772,16'd1359,-16'd2453,-16'd4586,-16'd7160,-16'd3936,-16'd2829,16'd645,-16'd4560,-16'd3214,16'd3150,-16'd6821,16'd2484,16'd2431,-16'd19,-16'd2514,-16'd4705,-16'd6722,-16'd5025,-16'd1705,-16'd760,16'd559,16'd4619,16'd4241,16'd775,16'd698,16'd4906,16'd7511,16'd6561,-16'd5380,16'd4898};
dout[292]={ -16'd49,-16'd7203,-16'd4244,16'd1661,-16'd5163,-16'd2417,-16'd4323,16'd4060,16'd5653,16'd9011,-16'd3908,-16'd7548,16'd2108,-16'd4968,16'd2970,16'd1963,-16'd39,-16'd1056,16'd4142,-16'd969,16'd3896,16'd2639,16'd2488,16'd3833,16'd172,-16'd6485,-16'd4612,16'd210,-16'd6786,-16'd5876,16'd1883,-16'd6286,-16'd2751,-16'd398,-16'd6960,16'd3702};
dout[293]={ 16'd288,16'd4542,-16'd3067,-16'd8386,16'd6672,16'd5238,-16'd332,16'd2120,16'd2510,-16'd4179,16'd6350,-16'd1762,-16'd4701,16'd5006,-16'd2908,16'd2192,16'd5659,16'd5757,-16'd165,-16'd5836,16'd9846,-16'd2340,16'd4192,-16'd3249,16'd8769,16'd2043,16'd135,16'd3494,16'd4249,16'd3941,-16'd4811,16'd416,16'd2384,16'd477,16'd2449,-16'd4929};
dout[294]={ -16'd964,16'd6110,-16'd5427,-16'd4331,16'd2888,-16'd1548,-16'd319,-16'd2270,16'd3745,-16'd529,16'd3077,-16'd2706,-16'd4420,-16'd228,16'd5102,16'd6936,-16'd2412,-16'd2030,-16'd3938,-16'd3878,-16'd3081,16'd5445,-16'd6646,-16'd7350,-16'd11,16'd5021,16'd4518,16'd5611,-16'd184,-16'd1780,-16'd34,-16'd499,-16'd8267,16'd4367,16'd4344,-16'd1052};
dout[295]={ -16'd5134,-16'd1309,16'd2397,16'd6586,-16'd6147,-16'd4286,-16'd1691,16'd580,16'd6445,16'd5736,-16'd6365,16'd440,16'd2577,-16'd5531,-16'd2923,-16'd7479,-16'd225,16'd4992,-16'd1056,16'd8038,16'd4222,-16'd6752,-16'd7438,16'd1190,-16'd320,16'd8599,-16'd7179,-16'd6791,-16'd199,16'd7834,-16'd4233,-16'd1973,16'd1287,16'd4361,16'd4538,16'd2078};
dout[296]={ -16'd5341,16'd3395,16'd3249,16'd3852,-16'd1321,-16'd7036,16'd4035,16'd1542,-16'd4127,-16'd1654,-16'd2204,16'd5668,16'd2317,16'd7322,16'd4,16'd2172,16'd7870,-16'd5052,-16'd6046,-16'd3264,-16'd5656,-16'd6907,16'd2958,16'd6456,-16'd2358,16'd6851,16'd2664,-16'd1392,16'd1048,16'd6951,16'd3819,-16'd6197,16'd4579,16'd5638,-16'd30,-16'd1515};
dout[297]={ 16'd4471,-16'd6316,-16'd1708,-16'd988,-16'd3122,-16'd4544,-16'd4525,-16'd5304,-16'd3410,-16'd2071,16'd3542,-16'd5895,-16'd3844,16'd5635,16'd3015,16'd6211,-16'd3936,-16'd4020,16'd7314,16'd4726,16'd3923,-16'd6867,-16'd6837,-16'd4273,-16'd380,-16'd1793,16'd1966,16'd2004,16'd112,16'd8058,16'd6932,-16'd5384,-16'd4080,-16'd1374,16'd4654,16'd10054};
dout[298]={ 16'd154,16'd4381,16'd7827,16'd3652,16'd1693,16'd1862,16'd1894,16'd2933,-16'd2639,-16'd3696,16'd388,16'd6118,-16'd5349,-16'd6738,16'd4245,-16'd3065,-16'd2248,16'd4989,-16'd7184,16'd2640,16'd3490,-16'd283,-16'd308,-16'd4748,16'd971,-16'd7251,-16'd6399,16'd2258,-16'd4644,16'd1618,-16'd5641,-16'd7226,16'd3753,-16'd5254,-16'd6780,16'd1518};
dout[299]={ 16'd3498,16'd5949,-16'd615,-16'd3483,16'd5378,16'd7421,16'd3659,16'd4896,-16'd5000,16'd7649,-16'd2151,-16'd3039,16'd439,16'd6578,-16'd6747,16'd630,-16'd1255,16'd5342,16'd6479,-16'd2792,16'd2002,16'd3221,-16'd6486,16'd7000,16'd1405,16'd2495,-16'd6706,-16'd4399,-16'd2690,16'd2964,-16'd5109,-16'd2188,-16'd136,16'd4445,16'd2186,16'd7000};
dout[300]={ 16'd8378,16'd5287,16'd5254,16'd6099,16'd227,16'd4574,-16'd2798,-16'd3435,16'd4163,16'd3885,-16'd12132,16'd3375,-16'd10448,-16'd588,16'd2767,16'd6393,16'd1790,-16'd4743,16'd5932,-16'd6628,16'd3079,-16'd4699,-16'd5441,-16'd87,16'd7273,16'd5584,16'd1872,-16'd5411,16'd5438,-16'd7538,-16'd4742,16'd3948,16'd348,16'd3995,16'd4351,-16'd923};
dout[301]={ 16'd2935,16'd9397,16'd2020,-16'd1338,-16'd2586,16'd8624,16'd6112,-16'd5270,16'd6551,16'd691,-16'd11265,-16'd6351,16'd1799,-16'd3920,-16'd4318,-16'd3822,16'd995,16'd1710,16'd432,-16'd2490,-16'd9443,16'd7,16'd8597,-16'd3922,16'd3385,16'd3137,16'd882,16'd802,16'd1458,16'd3172,-16'd5710,-16'd873,-16'd6406,-16'd4421,16'd5938,16'd3120};
dout[302]={ -16'd1019,16'd2034,-16'd3616,-16'd8543,16'd3216,-16'd6362,16'd4739,-16'd7415,16'd6155,-16'd3807,16'd4497,-16'd4004,16'd3173,-16'd8539,16'd2227,16'd1649,-16'd2821,16'd468,-16'd3609,-16'd5630,-16'd1487,-16'd3107,16'd2791,-16'd3709,16'd7036,-16'd5880,-16'd382,16'd3774,16'd2414,16'd6030,-16'd4860,16'd1809,16'd45,-16'd1424,-16'd2140,16'd7681};
dout[303]={ -16'd3443,-16'd382,16'd2188,16'd6035,16'd507,16'd2109,-16'd1547,-16'd2441,16'd6783,-16'd3233,-16'd5137,-16'd476,-16'd5716,16'd3106,-16'd983,16'd8829,-16'd9460,16'd5976,16'd4646,-16'd7046,-16'd2845,16'd3204,16'd6721,-16'd3345,-16'd3424,-16'd3806,-16'd4863,16'd1067,16'd438,-16'd1028,-16'd4129,16'd6592,-16'd3109,-16'd2708,-16'd3676,16'd357};
dout[304]={ -16'd4696,-16'd6686,16'd249,16'd5300,-16'd2157,16'd1513,16'd3054,-16'd8044,-16'd6039,-16'd1199,-16'd6679,-16'd1214,16'd2341,-16'd7579,-16'd4211,-16'd293,16'd4257,-16'd7841,16'd3627,16'd6131,-16'd3291,16'd1617,-16'd9628,16'd5795,16'd4674,-16'd4590,16'd871,-16'd3297,16'd3204,-16'd7483,16'd2307,-16'd6037,16'd4047,16'd3591,-16'd1665,-16'd4353};
dout[305]={ 16'd1457,-16'd1841,16'd5669,-16'd6926,16'd6217,-16'd2354,-16'd4322,-16'd22,-16'd393,16'd5952,-16'd1739,16'd5186,-16'd5563,16'd4770,16'd4978,16'd303,16'd6740,-16'd7378,-16'd6944,16'd6802,16'd1288,-16'd1418,16'd6133,16'd1134,-16'd1362,16'd2340,-16'd3783,-16'd45,16'd1339,-16'd7352,-16'd8226,-16'd713,16'd6187,-16'd6500,-16'd505,-16'd4501};
dout[306]={ 16'd2224,16'd6772,-16'd5224,16'd2204,16'd4303,-16'd4603,-16'd5050,16'd43,16'd3961,16'd4758,16'd4847,16'd3341,-16'd3940,16'd6546,-16'd499,16'd134,16'd790,-16'd6601,-16'd6075,-16'd3345,16'd5251,16'd2056,-16'd6559,16'd4892,16'd2102,16'd1182,-16'd3575,16'd7655,-16'd2936,-16'd4203,-16'd7108,-16'd4368,-16'd3927,-16'd3331,16'd3428,-16'd7569};
dout[307]={ -16'd4617,16'd4884,16'd6819,-16'd2097,16'd1699,16'd5402,16'd6832,-16'd7025,-16'd4702,-16'd3644,-16'd1006,16'd1463,16'd3337,-16'd3787,16'd4245,16'd4534,-16'd5535,-16'd1386,16'd6516,-16'd4053,-16'd6228,-16'd3248,16'd4944,-16'd5884,-16'd7781,-16'd1883,-16'd2137,16'd7573,16'd2471,16'd1752,-16'd1555,-16'd2370,-16'd3385,-16'd1117,-16'd5651,16'd5761};
dout[308]={ 16'd2291,16'd2904,-16'd2404,16'd861,16'd3106,16'd6685,-16'd3408,16'd6152,16'd4491,-16'd3491,-16'd1614,16'd2056,16'd3109,16'd2979,-16'd7214,-16'd4671,-16'd5206,-16'd2748,-16'd64,16'd3439,16'd7016,16'd1068,-16'd2523,-16'd6542,16'd735,-16'd205,16'd4202,-16'd6024,-16'd4048,16'd1809,-16'd5617,16'd1617,-16'd1626,-16'd7671,-16'd2234,-16'd4027};
dout[309]={ 16'd7469,-16'd2252,16'd723,16'd4852,16'd945,-16'd3505,16'd2763,-16'd1842,16'd2433,-16'd6445,16'd2027,-16'd2310,16'd1820,16'd1065,-16'd1571,-16'd969,-16'd2152,16'd4025,16'd5865,-16'd6542,-16'd1734,16'd5067,16'd4765,16'd3968,-16'd7617,16'd4585,16'd2983,16'd2952,-16'd6983,-16'd3525,16'd5838,-16'd4542,16'd1687,16'd7632,16'd6601,16'd2300};
dout[310]={ 16'd7311,-16'd3953,-16'd2654,-16'd2349,16'd5768,-16'd1850,-16'd7761,-16'd4847,16'd6516,16'd5198,-16'd8897,-16'd8315,-16'd7052,-16'd3671,16'd6375,16'd5799,-16'd5298,-16'd4359,16'd1696,16'd3889,16'd2820,16'd8244,-16'd748,-16'd5243,-16'd3636,16'd2007,16'd250,16'd4887,16'd2180,16'd1602,16'd8133,-16'd9460,-16'd1370,-16'd2033,16'd2705,-16'd27};
dout[311]={ 16'd2256,16'd3138,-16'd4969,16'd620,-16'd6507,16'd3383,-16'd137,16'd1778,16'd122,-16'd931,16'd748,-16'd1333,16'd5156,16'd330,16'd827,-16'd2982,-16'd4641,-16'd1702,16'd731,16'd2805,-16'd1631,-16'd4575,-16'd3268,16'd6564,16'd8554,-16'd2488,16'd3072,16'd184,-16'd5192,16'd9705,16'd1917,-16'd6772,-16'd2972,16'd694,-16'd4781,16'd6675};
dout[312]={ -16'd113,-16'd896,16'd1824,16'd1736,-16'd751,16'd3828,16'd5308,16'd92,-16'd5985,-16'd1102,-16'd6379,-16'd7086,16'd4079,-16'd6809,16'd1611,16'd5503,-16'd9427,-16'd6615,16'd7452,16'd2641,-16'd6895,-16'd792,16'd9176,-16'd5281,-16'd1675,-16'd1466,16'd4488,-16'd3719,-16'd742,16'd4990,16'd4391,-16'd4199,-16'd8258,16'd3144,-16'd5087,16'd7020};
dout[313]={ 16'd4270,-16'd6436,16'd1846,16'd1790,16'd1328,-16'd3221,-16'd574,16'd2284,16'd2165,16'd4760,16'd1832,16'd3618,16'd433,-16'd1784,16'd5642,16'd9025,-16'd3000,-16'd6556,-16'd1715,-16'd438,-16'd5477,-16'd2377,16'd1837,-16'd5815,-16'd5392,16'd5444,16'd4388,-16'd6319,-16'd4719,16'd3305,16'd8257,16'd6255,16'd517,-16'd935,-16'd5081,16'd5249};
dout[314]={ 16'd2247,16'd822,16'd55,16'd3935,16'd9001,16'd4824,-16'd1678,-16'd5498,16'd1186,16'd4041,16'd5034,-16'd6711,-16'd1726,-16'd1093,16'd5813,16'd617,16'd4605,16'd3561,16'd6637,16'd2248,16'd889,16'd8965,16'd2586,16'd4486,-16'd7845,16'd2487,16'd97,-16'd3521,-16'd4684,-16'd8443,-16'd4632,-16'd44,16'd4605,16'd3507,-16'd677,16'd5945};
dout[315]={ -16'd3880,-16'd2654,16'd6078,-16'd4612,16'd1167,-16'd5031,16'd2924,-16'd4165,16'd1028,-16'd3428,-16'd233,16'd4017,-16'd132,16'd4708,16'd84,-16'd4213,-16'd3936,-16'd4303,16'd5356,-16'd3574,-16'd362,16'd903,16'd441,16'd3371,16'd5230,-16'd2389,-16'd4945,16'd8133,-16'd3609,-16'd4591,16'd1523,-16'd6053,16'd4291,-16'd4135,16'd5268,-16'd4818};
dout[316]={ 16'd3803,-16'd845,-16'd1774,-16'd2826,16'd1323,-16'd6923,-16'd2361,-16'd1410,16'd2872,-16'd6634,-16'd4174,16'd5099,16'd177,-16'd7383,16'd1963,-16'd1183,-16'd1423,16'd3455,-16'd1520,16'd8042,16'd3964,16'd1888,16'd679,-16'd8965,-16'd4735,-16'd2312,-16'd4453,16'd2255,16'd5069,16'd1172,16'd3492,-16'd6868,16'd641,-16'd1918,-16'd7988,16'd5140};
dout[317]={ -16'd4401,-16'd2655,-16'd196,16'd2833,16'd4473,-16'd4862,16'd5582,16'd6131,-16'd2114,16'd4643,16'd2888,16'd5230,16'd5501,-16'd1134,-16'd2916,-16'd7110,16'd4608,-16'd609,16'd413,16'd5582,-16'd142,-16'd1484,16'd5631,16'd5804,16'd3240,16'd7385,16'd4289,16'd1573,16'd1396,-16'd2078,-16'd474,-16'd5047,-16'd2641,-16'd3785,16'd5197,-16'd2419};
dout[318]={ 16'd1079,-16'd2208,16'd8103,-16'd490,-16'd1113,16'd3926,-16'd2162,-16'd940,16'd449,-16'd678,-16'd4436,16'd5267,16'd3338,-16'd2274,-16'd3267,-16'd2570,16'd4935,16'd1614,-16'd3650,-16'd7507,16'd1822,16'd2641,16'd6288,16'd3139,-16'd129,16'd6377,16'd6793,-16'd835,-16'd4193,16'd6185,-16'd8140,16'd2353,16'd2229,-16'd5349,16'd820,-16'd2170};
dout[319]={ 16'd2299,16'd2663,16'd4414,-16'd6979,-16'd2408,16'd3511,-16'd3663,-16'd4499,16'd2203,-16'd4340,-16'd1569,-16'd3421,-16'd3804,16'd6382,16'd4354,16'd2142,-16'd5516,-16'd7577,16'd8013,-16'd5710,-16'd6298,16'd1636,-16'd5998,16'd4464,-16'd2255,-16'd8789,-16'd1225,16'd5399,16'd6189,16'd5541,-16'd3870,-16'd5491,16'd8105,-16'd2902,16'd736,16'd1140};
dout[320]={ -16'd4538,-16'd8116,-16'd2374,-16'd1043,-16'd4137,-16'd4678,-16'd179,16'd3867,-16'd5807,16'd2787,-16'd7500,16'd519,16'd830,-16'd6615,16'd2467,16'd11621,16'd5193,16'd1450,-16'd337,-16'd8784,-16'd1340,-16'd1923,-16'd8761,16'd2462,-16'd4665,-16'd1448,16'd3125,-16'd2564,-16'd399,16'd865,-16'd465,16'd571,-16'd13108,16'd3686,-16'd3062,16'd5112};
dout[321]={ 16'd4583,16'd3864,-16'd2974,-16'd1280,16'd8039,16'd2934,16'd7842,-16'd414,-16'd3838,-16'd5688,-16'd4770,16'd796,16'd4192,-16'd478,16'd6923,-16'd4308,16'd2055,-16'd5734,16'd5008,16'd3872,16'd3183,-16'd5769,16'd6312,-16'd4935,16'd9329,-16'd2464,-16'd1297,-16'd9207,-16'd6832,16'd7449,-16'd369,-16'd2690,-16'd2262,16'd1653,16'd5196,-16'd2389};
dout[322]={ 16'd1239,16'd6408,-16'd7928,16'd2357,-16'd5643,-16'd3970,-16'd1703,16'd3088,-16'd602,-16'd3472,-16'd5910,-16'd4412,16'd1899,-16'd1565,16'd1211,16'd3297,-16'd4410,16'd7774,16'd5563,-16'd2831,-16'd2949,-16'd7153,16'd8388,16'd4917,16'd3280,-16'd2911,16'd266,16'd550,16'd991,16'd10161,16'd9034,-16'd1126,-16'd351,-16'd2705,16'd2240,16'd6083};
dout[323]={ -16'd4210,16'd8464,-16'd4573,-16'd3102,-16'd991,16'd3055,-16'd305,16'd4475,-16'd7605,-16'd5994,-16'd8176,-16'd3166,-16'd3929,-16'd6937,16'd2084,16'd265,-16'd4059,-16'd3239,-16'd6189,-16'd5291,16'd6785,-16'd1040,-16'd5575,-16'd6466,-16'd2376,-16'd8695,-16'd4147,16'd4353,-16'd2031,-16'd3613,-16'd3737,16'd1095,-16'd10378,16'd4132,-16'd5997,-16'd4742};
dout[324]={ 16'd8484,-16'd7072,-16'd3800,16'd4104,16'd5009,16'd3219,-16'd2857,16'd3739,-16'd4227,-16'd572,-16'd4035,-16'd4426,16'd1266,-16'd4552,-16'd6116,16'd2575,-16'd655,-16'd5303,16'd4991,16'd1712,16'd5350,16'd3233,-16'd7747,16'd3536,-16'd1781,16'd3894,-16'd1419,16'd3772,16'd2710,16'd4735,-16'd5201,16'd5028,16'd4077,16'd4352,-16'd7094,-16'd6140};
dout[325]={ 16'd1602,16'd5273,-16'd1416,-16'd3245,16'd6250,16'd1573,16'd24,16'd1996,-16'd3772,-16'd4907,16'd4338,16'd1744,16'd4052,-16'd6207,-16'd3608,-16'd7764,16'd3870,-16'd3119,-16'd2294,16'd1208,16'd4071,-16'd1318,16'd1954,-16'd4728,16'd2092,-16'd4550,-16'd2992,16'd2574,-16'd8107,-16'd2914,-16'd2330,16'd5219,-16'd4843,16'd1901,-16'd790,-16'd1796};
dout[326]={ -16'd3779,-16'd4203,-16'd5555,-16'd7182,-16'd3083,16'd5663,16'd585,16'd6618,16'd4768,16'd5117,-16'd862,16'd1504,-16'd1594,-16'd1589,-16'd4743,16'd249,-16'd5689,-16'd5904,-16'd7221,-16'd6517,16'd2770,16'd4456,-16'd2059,16'd4830,-16'd1824,-16'd989,-16'd4288,-16'd4392,-16'd5243,-16'd2835,16'd7609,16'd2427,-16'd3958,-16'd868,-16'd5967,16'd2808};
dout[327]={ -16'd1037,16'd420,16'd3461,-16'd7272,16'd1686,-16'd6106,-16'd4370,-16'd90,16'd2833,16'd2525,-16'd2908,16'd3792,-16'd4077,-16'd5101,16'd2242,-16'd2719,16'd4837,16'd307,16'd151,16'd1787,-16'd4330,-16'd7439,16'd1591,16'd5313,-16'd610,-16'd3938,-16'd4966,16'd814,16'd4603,-16'd6723,-16'd5553,-16'd5384,16'd1428,-16'd3897,16'd6007,16'd3828};
dout[328]={ -16'd6376,-16'd1995,16'd5961,16'd5558,16'd4299,16'd2988,-16'd4258,16'd3857,16'd2013,16'd3441,-16'd2809,16'd4609,16'd4004,16'd3466,-16'd4060,-16'd2689,-16'd2563,-16'd2581,-16'd3580,16'd1191,-16'd5722,16'd680,-16'd4002,-16'd4532,-16'd6239,16'd4475,-16'd3087,16'd2735,-16'd7474,-16'd5674,16'd5162,-16'd6766,-16'd1270,-16'd6213,16'd889,16'd5915};
dout[329]={ 16'd2070,-16'd173,16'd730,-16'd8319,-16'd3661,-16'd4887,16'd5678,-16'd3953,-16'd4120,16'd2383,16'd767,-16'd6169,-16'd4614,16'd5068,16'd3525,16'd1541,16'd6007,-16'd6379,16'd8480,16'd5995,-16'd6438,16'd4784,16'd132,-16'd3199,16'd3176,-16'd3508,16'd3869,16'd451,-16'd3262,16'd6302,16'd7992,16'd526,-16'd2061,16'd3234,16'd4134,-16'd6436};
dout[330]={ -16'd57,16'd912,-16'd5548,-16'd3503,16'd3406,-16'd8004,16'd7110,16'd399,-16'd9562,-16'd5570,16'd3558,16'd1458,16'd714,-16'd90,-16'd809,16'd3524,16'd740,-16'd8343,16'd1966,-16'd4141,16'd839,-16'd3164,-16'd3913,-16'd5857,-16'd3352,-16'd2902,16'd2041,-16'd4690,16'd4793,16'd4673,-16'd147,-16'd4633,-16'd8195,16'd4618,16'd1801,-16'd5792};
dout[331]={ 16'd2121,-16'd3849,-16'd102,-16'd522,16'd2127,-16'd5350,-16'd6537,16'd6499,16'd404,16'd6436,-16'd11295,-16'd7446,16'd2975,-16'd1704,-16'd8315,-16'd1304,-16'd6428,16'd7020,16'd3318,-16'd2119,16'd7333,16'd7722,16'd4920,-16'd6416,16'd8501,-16'd2132,-16'd7072,16'd4729,16'd2758,16'd4202,16'd10519,16'd4480,-16'd12264,-16'd1213,-16'd4584,16'd2638};
dout[332]={ -16'd2174,-16'd4808,-16'd5912,16'd743,-16'd6375,-16'd1301,-16'd451,-16'd280,-16'd4976,16'd4296,-16'd13968,-16'd2627,16'd4441,-16'd9220,-16'd2682,16'd4516,-16'd2369,16'd598,-16'd1143,-16'd2982,16'd886,16'd6858,16'd5336,-16'd6504,16'd4082,-16'd73,-16'd4405,16'd158,16'd689,16'd8631,16'd5606,16'd2699,-16'd13050,-16'd5061,16'd1370,16'd1680};
dout[333]={ 16'd5976,16'd1267,16'd5261,16'd2213,-16'd2082,-16'd3048,-16'd6392,16'd342,16'd6608,16'd5155,-16'd7449,16'd5674,-16'd6856,16'd4410,-16'd979,-16'd906,16'd4473,16'd913,16'd1056,16'd4169,16'd435,-16'd3480,16'd5886,-16'd7925,16'd6155,-16'd1189,-16'd2753,16'd3234,16'd4869,-16'd3439,16'd8985,16'd1396,-16'd5046,-16'd8506,-16'd8869,16'd5590};
dout[334]={ -16'd2221,16'd1650,16'd1532,16'd1277,-16'd199,16'd6677,16'd8546,-16'd6369,16'd4068,-16'd620,16'd5701,-16'd5226,-16'd4106,16'd2257,-16'd1191,16'd4776,16'd665,-16'd5300,-16'd7994,-16'd7107,16'd607,16'd6959,-16'd7919,16'd4989,16'd3614,-16'd1630,-16'd369,16'd6758,-16'd5078,-16'd2044,16'd6731,-16'd2719,-16'd5000,16'd512,16'd490,-16'd5435};
dout[335]={ -16'd111,-16'd6683,-16'd8787,-16'd6235,-16'd4428,-16'd6562,16'd8051,16'd2768,16'd2670,-16'd4276,16'd8145,16'd304,16'd28,16'd5933,16'd647,-16'd427,16'd4891,16'd659,16'd2224,-16'd2189,-16'd6616,16'd936,16'd7998,-16'd1793,-16'd289,16'd3981,16'd6694,16'd2142,-16'd6841,16'd5295,16'd5484,16'd1267,-16'd264,-16'd1954,16'd537,16'd883};
dout[336]={ 16'd3675,16'd3245,16'd1264,16'd2903,16'd791,-16'd3141,-16'd1076,16'd2497,-16'd1772,16'd3002,-16'd1522,16'd5865,-16'd405,16'd3469,-16'd4858,-16'd5310,-16'd384,-16'd3445,-16'd7027,16'd5207,16'd7212,16'd1691,-16'd1447,16'd2826,-16'd3832,16'd7278,-16'd5745,16'd4948,16'd4961,-16'd2273,16'd6267,-16'd1738,-16'd2578,-16'd3273,16'd4704,16'd343};
dout[337]={ -16'd2334,16'd6064,16'd2791,-16'd3043,16'd6172,16'd269,-16'd2611,-16'd3033,-16'd2893,16'd3485,16'd2685,16'd278,-16'd2858,16'd6983,-16'd1274,16'd4096,-16'd4264,16'd4108,16'd5203,16'd12,16'd4278,-16'd6168,16'd1074,-16'd5166,-16'd839,-16'd1113,-16'd3101,16'd2568,16'd1780,16'd4558,-16'd1084,-16'd439,16'd1054,-16'd6466,-16'd4144,-16'd1171};
dout[338]={ -16'd2437,-16'd1394,-16'd1024,-16'd2401,16'd7910,-16'd844,-16'd4503,-16'd2240,-16'd2475,-16'd7246,-16'd2484,16'd1201,-16'd391,16'd3917,-16'd5360,16'd3099,16'd7192,16'd7070,-16'd5986,-16'd4720,16'd6949,-16'd4974,-16'd2648,-16'd3424,16'd1771,16'd1140,-16'd6778,-16'd396,16'd2650,16'd593,16'd5811,-16'd6542,-16'd6439,16'd2244,16'd3599,16'd1272};
dout[339]={ -16'd5304,-16'd73,-16'd8834,16'd624,16'd190,16'd2011,16'd5730,16'd7009,-16'd6393,16'd5583,16'd7385,16'd16,16'd3258,-16'd4276,16'd2867,-16'd3985,-16'd5686,-16'd4930,16'd8143,16'd8821,16'd1899,16'd1676,-16'd5352,-16'd3424,-16'd3185,16'd763,16'd4481,16'd5717,16'd5614,-16'd372,-16'd502,16'd734,-16'd4301,16'd3542,-16'd7466,-16'd2911};
dout[340]={ -16'd8505,-16'd3667,-16'd4683,16'd3204,-16'd235,-16'd13527,-16'd281,-16'd4915,-16'd9762,16'd8911,16'd3125,-16'd54,-16'd2291,16'd3658,-16'd9332,16'd5125,-16'd3172,-16'd4033,16'd5704,-16'd9418,16'd1310,-16'd2763,-16'd8811,-16'd1323,-16'd3534,16'd5035,-16'd219,16'd2273,-16'd3653,16'd1229,16'd6622,16'd1913,-16'd16714,16'd4797,-16'd108,16'd5758};
dout[341]={ 16'd4905,-16'd6964,16'd3285,16'd2840,-16'd4903,16'd2659,16'd1073,-16'd2535,-16'd4714,16'd2651,-16'd9977,-16'd3624,16'd2796,16'd5824,-16'd7541,-16'd4266,16'd6058,16'd9272,16'd7833,-16'd7716,16'd7977,16'd2380,-16'd1008,-16'd6175,16'd5809,-16'd6728,-16'd6066,-16'd1077,16'd3305,16'd2323,16'd3311,-16'd695,-16'd2674,16'd3273,16'd132,-16'd2682};
dout[342]={ -16'd7938,-16'd6584,16'd3382,-16'd4042,-16'd864,-16'd2270,-16'd5017,-16'd3021,16'd4705,16'd5552,-16'd5428,-16'd7482,-16'd1187,16'd3045,-16'd8471,16'd5638,-16'd6460,16'd2687,16'd4620,-16'd6930,-16'd6666,-16'd9741,-16'd1402,-16'd392,16'd9566,-16'd7690,-16'd3271,16'd3483,16'd4184,-16'd2545,16'd6924,-16'd7496,-16'd7273,16'd8878,16'd1813,16'd6980};
dout[343]={ 16'd3299,-16'd4068,-16'd8713,16'd3423,-16'd8732,16'd346,-16'd5395,-16'd7602,-16'd4740,16'd8629,-16'd1327,16'd4974,16'd4404,16'd5774,-16'd8882,16'd146,16'd662,-16'd4575,16'd2998,-16'd3780,16'd7382,16'd3480,-16'd4005,-16'd9428,-16'd1807,-16'd6980,16'd6757,-16'd362,-16'd4692,-16'd837,16'd5683,-16'd5772,16'd5040,-16'd701,16'd2559,-16'd1605};
dout[344]={ -16'd2271,16'd5784,16'd244,16'd6211,16'd6467,-16'd5767,-16'd7941,16'd3255,-16'd584,-16'd7492,16'd3619,-16'd3183,16'd2666,-16'd1354,-16'd7772,-16'd5805,16'd1825,16'd566,-16'd8842,-16'd7993,-16'd207,16'd2264,-16'd6830,16'd680,16'd2624,-16'd6430,-16'd54,-16'd4552,-16'd1800,-16'd7160,-16'd451,-16'd761,16'd459,16'd511,-16'd2420,-16'd4728};
dout[345]={ -16'd3774,16'd4035,-16'd2836,16'd1896,-16'd2848,16'd2340,16'd6791,16'd2531,16'd890,16'd6635,16'd4405,16'd4347,16'd5493,16'd2142,16'd5765,16'd292,16'd6177,-16'd4432,16'd5333,-16'd5786,-16'd3801,16'd7791,-16'd4841,-16'd235,-16'd2886,-16'd1003,-16'd580,-16'd3529,-16'd633,-16'd3561,16'd7489,-16'd4216,-16'd6731,-16'd647,16'd3452,16'd505};
dout[346]={ 16'd5316,16'd3662,-16'd2220,16'd2673,-16'd3770,-16'd6346,16'd2156,-16'd570,-16'd1849,-16'd4570,-16'd3336,16'd2114,-16'd7307,16'd3682,-16'd2013,16'd1062,-16'd6245,-16'd3669,-16'd6930,16'd2642,-16'd5988,-16'd6363,16'd2034,-16'd3534,16'd4589,16'd1392,16'd4011,16'd1449,16'd4573,16'd6303,-16'd2573,-16'd1438,-16'd4321,-16'd5902,16'd1990,16'd1088};
dout[347]={ 16'd5873,16'd2906,16'd5845,-16'd9318,16'd4360,16'd6055,-16'd2722,-16'd6390,-16'd2910,16'd636,16'd4469,-16'd5008,16'd2389,-16'd3710,-16'd6849,-16'd4122,16'd2774,-16'd4882,-16'd6457,16'd5616,-16'd4683,16'd5185,-16'd1502,-16'd112,-16'd2688,-16'd3247,-16'd2963,-16'd3680,16'd4782,16'd3751,16'd6100,-16'd751,16'd2863,-16'd1425,16'd6466,16'd4545};
dout[348]={ 16'd3958,-16'd1924,-16'd8239,16'd2465,16'd2975,16'd2151,-16'd5542,-16'd9082,16'd499,16'd1040,-16'd4467,-16'd338,-16'd6375,16'd4678,-16'd2014,-16'd779,-16'd1002,16'd8101,-16'd4944,16'd2492,16'd6059,-16'd5151,-16'd2590,16'd6784,16'd514,16'd482,16'd1447,16'd2124,16'd3197,-16'd6283,-16'd7999,16'd4957,16'd6806,16'd5393,-16'd6945,16'd6336};
dout[349]={ 16'd6548,16'd3639,-16'd2014,-16'd509,16'd8799,-16'd4446,-16'd1382,16'd6843,16'd3311,16'd4685,16'd6661,-16'd2535,16'd1902,16'd3626,16'd763,16'd2580,-16'd3274,-16'd2728,16'd818,16'd2460,-16'd6408,-16'd3267,16'd5885,16'd7236,16'd4389,16'd5690,-16'd4565,16'd3100,-16'd5099,16'd4637,-16'd5995,16'd3322,-16'd745,-16'd718,16'd1413,16'd1824};
dout[350]={ -16'd7276,-16'd762,16'd4315,16'd912,-16'd6678,-16'd11357,16'd2532,-16'd4704,-16'd6157,16'd4415,16'd568,-16'd8724,16'd478,16'd7601,-16'd1723,16'd8803,-16'd373,-16'd6203,16'd4047,-16'd5448,-16'd7076,16'd3078,-16'd1452,16'd411,16'd3626,16'd10379,-16'd3917,-16'd4185,16'd2790,-16'd1198,-16'd2169,16'd1396,-16'd13836,-16'd3361,-16'd1581,-16'd5152};
dout[351]={ -16'd7115,-16'd545,-16'd4201,-16'd6521,-16'd4983,16'd556,-16'd6212,-16'd5721,-16'd931,-16'd4294,-16'd1164,-16'd4700,16'd1143,16'd2618,16'd5606,-16'd2187,-16'd1643,16'd5974,-16'd1611,-16'd4378,16'd2658,-16'd8952,-16'd5873,-16'd1063,16'd3889,-16'd9920,-16'd5611,16'd5916,16'd6406,16'd4546,-16'd4794,16'd928,-16'd354,16'd8974,-16'd8807,-16'd6837};
dout[352]={ -16'd10432,16'd489,-16'd4436,-16'd961,-16'd2176,-16'd10822,-16'd8194,16'd8376,-16'd498,-16'd5144,-16'd2366,-16'd10266,16'd4896,-16'd2824,16'd4045,16'd591,-16'd599,16'd8268,16'd512,-16'd3011,-16'd2920,-16'd6677,16'd1861,-16'd6430,-16'd3912,-16'd9029,-16'd7182,-16'd5314,-16'd3917,-16'd5714,-16'd1909,16'd639,16'd2909,-16'd4874,-16'd4881,-16'd7819};
dout[353]={ 16'd7366,-16'd1701,-16'd3336,-16'd3560,16'd3749,16'd1536,16'd5220,16'd1641,-16'd3179,16'd6084,16'd2679,-16'd7294,16'd3169,-16'd3404,-16'd5005,-16'd2962,16'd1543,16'd1652,-16'd7352,-16'd8574,16'd6890,-16'd7434,16'd7167,-16'd3315,-16'd4926,-16'd1224,-16'd6790,-16'd1491,16'd3105,-16'd8847,-16'd4036,-16'd5644,16'd1159,16'd4511,16'd4856,-16'd180};
dout[354]={ 16'd9841,-16'd5287,-16'd5734,16'd4981,-16'd5598,-16'd1982,16'd2931,-16'd4821,-16'd3290,-16'd5,16'd4899,16'd3679,16'd5464,-16'd4043,-16'd7085,16'd3604,16'd3660,-16'd7657,16'd4439,16'd2433,16'd1498,16'd3334,16'd1471,-16'd6476,-16'd3015,-16'd7171,16'd1406,-16'd509,16'd3636,16'd5374,16'd6558,16'd4706,-16'd3291,-16'd616,-16'd864,16'd12};
dout[355]={ 16'd138,16'd1488,-16'd1940,-16'd2860,16'd2002,-16'd2511,16'd715,-16'd4976,16'd2307,16'd3254,16'd3103,16'd3488,16'd1502,16'd388,16'd5272,-16'd4815,-16'd1362,16'd3855,-16'd5754,16'd5192,16'd3663,16'd755,-16'd2088,-16'd4416,16'd5284,-16'd815,16'd2385,16'd2488,16'd1515,-16'd1027,16'd2481,-16'd4065,-16'd2860,-16'd1068,-16'd43,16'd5883};
dout[356]={ 16'd6466,16'd3147,16'd6431,16'd3641,16'd2106,-16'd4798,-16'd258,16'd1486,16'd6134,16'd6714,16'd5504,16'd332,16'd3539,16'd7312,16'd2026,16'd369,16'd3932,-16'd6414,16'd6226,16'd3136,16'd2239,16'd1548,-16'd2403,-16'd246,16'd7711,-16'd1850,-16'd2911,16'd3980,16'd5175,-16'd4614,16'd3427,-16'd3135,-16'd3931,16'd1570,-16'd3509,16'd5721};
dout[357]={ -16'd1450,16'd746,16'd5336,-16'd6206,16'd1191,16'd6174,16'd3889,16'd5133,-16'd1657,16'd3830,16'd1887,-16'd4749,-16'd772,-16'd3699,16'd5489,16'd1997,16'd4855,-16'd1887,16'd1381,16'd5932,-16'd4962,16'd4819,16'd5036,16'd7125,16'd4182,-16'd397,-16'd6126,16'd5590,16'd3280,16'd5558,16'd1973,-16'd734,16'd2862,16'd4648,-16'd4740,16'd4486};
dout[358]={ -16'd3200,-16'd4049,16'd1035,16'd1138,-16'd1382,16'd265,-16'd5947,-16'd7957,-16'd3400,16'd2568,-16'd2955,-16'd2899,-16'd3571,16'd7338,16'd123,16'd5864,-16'd4559,16'd5861,16'd4306,16'd7140,-16'd2065,-16'd1264,-16'd635,-16'd4808,16'd5355,16'd884,16'd2847,16'd1217,16'd2939,-16'd3042,16'd1824,-16'd1654,16'd3909,-16'd850,-16'd2243,-16'd5049};
dout[359]={ 16'd797,16'd7717,16'd5622,-16'd335,16'd2972,16'd4760,16'd4980,-16'd2037,-16'd6182,16'd7518,16'd5418,16'd4223,16'd5698,16'd6935,-16'd2340,-16'd1020,-16'd4272,16'd7305,16'd1554,-16'd146,16'd5204,16'd2975,-16'd7379,16'd5203,16'd2367,-16'd3361,16'd6227,16'd4231,16'd1182,16'd7330,16'd4597,16'd1613,16'd2875,-16'd3621,16'd6828,16'd5022};
dout[360]={ 16'd406,-16'd3221,16'd2752,16'd658,-16'd1073,-16'd8080,-16'd5103,16'd2715,16'd2887,16'd10939,16'd3260,16'd468,-16'd2190,-16'd3308,-16'd3981,16'd5313,-16'd3086,-16'd8343,-16'd2052,16'd884,-16'd8885,-16'd409,-16'd7447,-16'd1027,16'd4076,16'd5595,16'd7336,16'd5925,16'd4494,-16'd2804,16'd3833,-16'd2715,-16'd2503,16'd4990,-16'd5027,-16'd6583};
dout[361]={ -16'd3991,-16'd6012,-16'd3148,-16'd6620,-16'd5948,-16'd8089,-16'd4978,-16'd2016,-16'd6577,16'd2249,-16'd4894,16'd5182,16'd3702,16'd10135,-16'd8,-16'd3354,-16'd1682,16'd659,16'd3166,-16'd7091,16'd862,-16'd8237,-16'd6993,-16'd6244,16'd6643,16'd450,-16'd270,16'd605,-16'd2271,-16'd2904,-16'd6410,-16'd7960,16'd3159,-16'd4563,-16'd9251,16'd6064};
dout[362]={ -16'd6227,-16'd7871,-16'd4600,-16'd2553,-16'd62,-16'd3886,16'd2001,-16'd4940,16'd1499,-16'd6331,-16'd8119,-16'd3234,16'd5103,-16'd219,16'd5468,16'd684,-16'd4351,16'd4220,-16'd7958,-16'd175,-16'd5479,-16'd2073,-16'd409,-16'd3454,16'd3325,-16'd9548,-16'd5991,-16'd1289,-16'd422,-16'd2861,-16'd1769,-16'd1634,-16'd1734,16'd6139,16'd1948,16'd230};
dout[363]={ 16'd500,16'd6239,16'd7821,16'd739,-16'd6322,-16'd12385,16'd1996,-16'd7711,-16'd8607,-16'd5274,16'd445,16'd2233,16'd1538,16'd3685,16'd3692,16'd3816,16'd8253,-16'd1645,-16'd8396,-16'd9264,16'd3441,16'd1411,-16'd3129,-16'd8057,16'd4855,16'd4022,-16'd686,16'd2598,-16'd1506,16'd5357,16'd6680,16'd2514,16'd4107,-16'd1101,-16'd1746,16'd7394};
dout[364]={ 16'd7571,16'd631,-16'd5209,16'd7100,-16'd2539,-16'd5313,-16'd297,16'd8505,-16'd1187,16'd3093,16'd9490,16'd5995,16'd3839,16'd3886,-16'd9674,16'd1416,-16'd3192,-16'd8837,-16'd9134,-16'd4435,-16'd2322,-16'd8372,16'd1831,16'd4606,-16'd1764,-16'd2729,-16'd4116,-16'd5345,-16'd4404,-16'd4840,-16'd6256,-16'd4466,16'd2839,-16'd6309,-16'd965,-16'd5015};
dout[365]={ 16'd4323,-16'd6110,-16'd3822,16'd8437,16'd5586,16'd3035,-16'd5648,-16'd276,-16'd7120,16'd2603,16'd8037,-16'd1905,16'd4328,16'd3204,16'd4160,-16'd6979,-16'd6203,-16'd1737,-16'd1019,16'd1143,-16'd2051,16'd4079,16'd5760,16'd1639,16'd715,-16'd1878,16'd1663,-16'd797,16'd4212,16'd6750,-16'd4118,-16'd2460,16'd1990,16'd4541,16'd534,-16'd5359};
dout[366]={ 16'd3170,-16'd4669,16'd4444,-16'd4448,-16'd2653,16'd1438,-16'd5020,-16'd2433,-16'd4251,-16'd5757,-16'd4177,-16'd3710,-16'd5359,-16'd2094,-16'd1179,16'd5560,-16'd613,-16'd8356,-16'd3180,-16'd1772,-16'd1165,-16'd7068,-16'd4608,-16'd5497,-16'd3039,16'd6329,16'd3464,16'd2610,-16'd3633,16'd5655,-16'd3398,16'd2584,16'd479,-16'd6474,-16'd5356,16'd3195};
dout[367]={ -16'd1544,-16'd1740,16'd162,16'd1576,-16'd1283,16'd564,-16'd2296,16'd1661,16'd4652,16'd1552,16'd3849,16'd750,16'd5595,-16'd2726,16'd3787,16'd3675,16'd4034,-16'd6108,-16'd6179,-16'd1386,16'd235,-16'd7427,16'd4544,16'd4064,-16'd3231,16'd5270,-16'd197,-16'd5979,16'd3645,16'd6946,-16'd3624,-16'd5939,16'd6163,-16'd999,16'd4304,16'd4450};
dout[368]={ 16'd4331,16'd2399,-16'd8290,16'd1749,16'd4081,-16'd4881,-16'd6040,-16'd4114,16'd4973,16'd3397,16'd5584,-16'd4994,16'd4595,-16'd1307,-16'd1998,-16'd1678,-16'd3271,16'd4583,16'd858,-16'd2403,-16'd448,-16'd6403,16'd2484,16'd2251,-16'd5601,16'd6273,-16'd2165,-16'd3317,-16'd6204,16'd2571,16'd5672,-16'd2173,16'd7110,16'd4273,-16'd4542,16'd5377};
dout[369]={ -16'd3787,16'd7584,16'd756,-16'd3547,16'd4977,-16'd4430,-16'd5063,-16'd6942,-16'd783,-16'd3158,-16'd2042,16'd8081,16'd23,-16'd929,-16'd3383,-16'd4720,16'd3510,-16'd487,16'd6163,-16'd2745,16'd6024,16'd3372,-16'd258,-16'd290,-16'd988,-16'd6492,-16'd4418,-16'd5460,-16'd969,16'd1186,16'd3122,-16'd7317,-16'd6094,16'd224,16'd7005,16'd3820};
dout[370]={ 16'd347,-16'd12437,16'd2380,16'd603,-16'd5157,-16'd642,16'd512,16'd714,-16'd8064,16'd6275,16'd539,-16'd4823,-16'd235,16'd3712,16'd1620,16'd11375,16'd774,-16'd6491,-16'd1069,16'd307,-16'd6666,16'd123,16'd548,16'd172,16'd4449,16'd1469,16'd8631,16'd2408,16'd978,-16'd3448,16'd2696,-16'd9024,16'd4639,-16'd1557,-16'd4015,-16'd190};
dout[371]={ -16'd4949,-16'd6207,-16'd1827,-16'd2167,-16'd7775,16'd4148,16'd793,16'd1114,-16'd3404,-16'd1315,-16'd3140,-16'd7156,-16'd6597,16'd2570,-16'd6275,-16'd4491,16'd1581,-16'd2210,-16'd664,-16'd5591,16'd3149,-16'd4772,-16'd1281,-16'd8365,-16'd1736,16'd5286,-16'd5326,-16'd95,-16'd4755,-16'd774,-16'd8574,-16'd8744,16'd4570,-16'd1010,-16'd5760,16'd380};
dout[372]={ -16'd98,16'd1827,-16'd5025,-16'd8300,16'd1177,-16'd8454,-16'd4014,-16'd3430,-16'd6568,-16'd6533,-16'd3183,16'd2806,16'd2402,16'd4995,-16'd9576,-16'd1388,-16'd1345,16'd4290,-16'd571,16'd3932,-16'd3010,-16'd7507,16'd4788,-16'd4767,-16'd2599,-16'd4509,16'd5421,16'd8546,-16'd4711,16'd836,-16'd8254,16'd1792,-16'd10606,-16'd2525,16'd437,16'd5105};
dout[373]={ -16'd1503,-16'd7041,-16'd2570,-16'd3422,-16'd5494,-16'd13092,16'd2986,-16'd213,16'd2470,16'd4063,16'd10803,-16'd7600,16'd2664,-16'd2087,-16'd7073,-16'd1166,16'd10591,16'd211,-16'd8482,-16'd3831,-16'd4989,-16'd2658,16'd2214,-16'd3881,-16'd7648,16'd5451,-16'd7618,-16'd2029,-16'd1708,-16'd3918,-16'd6390,16'd4229,16'd1522,16'd2827,-16'd613,16'd7820};
dout[374]={ 16'd7077,-16'd4628,-16'd3570,16'd12951,-16'd6041,16'd6165,16'd7200,16'd2306,16'd2240,-16'd337,-16'd2030,-16'd3525,-16'd6510,16'd4727,16'd2341,-16'd551,16'd6967,16'd3004,16'd3792,-16'd3547,-16'd6131,16'd4848,-16'd6770,-16'd3763,16'd4293,16'd6510,16'd129,-16'd7258,16'd4640,16'd1257,-16'd3312,-16'd1719,16'd8945,16'd6576,16'd7936,-16'd2589};
dout[375]={ -16'd2610,-16'd6909,16'd376,16'd3016,-16'd6344,16'd5940,16'd6550,-16'd3231,-16'd4266,16'd4113,-16'd5051,-16'd3337,16'd7998,16'd2054,-16'd7798,16'd981,16'd437,-16'd3759,-16'd7104,16'd1542,-16'd1743,-16'd3211,-16'd3821,16'd1291,-16'd212,-16'd1887,16'd2321,16'd292,16'd2124,-16'd3887,-16'd5684,-16'd7023,-16'd2990,16'd4894,-16'd4173,-16'd4658};
dout[376]={ 16'd3763,16'd7684,-16'd2276,-16'd2483,-16'd1577,16'd7457,16'd5904,-16'd3347,-16'd4968,-16'd1515,16'd4484,16'd993,-16'd4621,-16'd4361,16'd5958,-16'd5748,-16'd6041,-16'd1342,16'd451,16'd3944,-16'd162,16'd2284,16'd2202,16'd4945,16'd6553,16'd270,-16'd1559,-16'd5461,16'd6324,16'd852,-16'd160,-16'd7557,16'd5197,16'd1779,-16'd1350,-16'd7568};
dout[377]={ -16'd1412,-16'd2344,-16'd4162,16'd1301,-16'd2978,16'd500,-16'd6304,-16'd5194,-16'd3024,-16'd6409,16'd4024,-16'd6058,16'd3405,-16'd3748,16'd5127,16'd2960,16'd4921,16'd6141,-16'd6183,-16'd3049,16'd4300,16'd4509,-16'd4278,16'd6701,16'd6631,16'd4959,-16'd1550,16'd4554,16'd5480,-16'd735,-16'd4786,16'd3263,-16'd3274,16'd5427,16'd6502,-16'd4012};
dout[378]={ -16'd8570,-16'd5590,16'd1299,16'd3029,-16'd5146,-16'd3047,16'd55,-16'd4602,16'd2803,16'd770,16'd3204,16'd3511,-16'd5248,16'd109,16'd8993,-16'd4254,-16'd3905,16'd1513,16'd6120,-16'd166,16'd2362,-16'd570,-16'd1795,16'd2870,-16'd4780,-16'd246,-16'd3233,16'd6314,16'd2650,16'd79,-16'd2991,16'd1593,16'd466,16'd6127,-16'd4017,16'd1087};
dout[379]={ -16'd7747,16'd299,-16'd4417,16'd2946,16'd1309,-16'd403,16'd4445,-16'd7202,-16'd5175,16'd94,-16'd274,-16'd729,-16'd1859,-16'd4166,16'd3961,16'd4214,16'd4179,16'd5874,-16'd5368,16'd2775,16'd3227,16'd3271,-16'd7299,-16'd6651,16'd3823,-16'd1256,16'd1717,16'd3492,16'd372,16'd1973,16'd2216,-16'd7510,-16'd2152,-16'd5161,-16'd4822,-16'd7479};
dout[380]={ -16'd8374,-16'd16707,-16'd4036,16'd3223,-16'd1076,16'd4180,-16'd793,16'd3077,16'd4594,-16'd2764,-16'd5911,16'd2586,16'd2442,-16'd8940,-16'd6932,16'd8207,16'd1136,-16'd10001,16'd3350,-16'd2734,16'd5573,-16'd802,16'd251,-16'd4565,16'd3118,16'd10393,16'd7017,16'd4970,-16'd1025,-16'd4713,-16'd6436,-16'd5240,16'd8257,16'd3514,-16'd5314,-16'd8791};
dout[381]={ 16'd3330,-16'd7592,16'd5799,-16'd5949,-16'd6281,-16'd627,16'd1592,-16'd887,16'd1481,-16'd8012,16'd4116,16'd2874,16'd3693,16'd249,-16'd3781,-16'd1433,-16'd4454,16'd2985,-16'd2555,-16'd6514,-16'd7998,-16'd2081,16'd1154,16'd4468,-16'd1032,16'd4481,-16'd6880,16'd8169,-16'd9099,16'd5581,-16'd1312,16'd1921,-16'd1879,-16'd8765,-16'd5612,-16'd2791};
dout[382]={ -16'd6527,16'd1629,16'd5119,-16'd9707,-16'd11693,-16'd12362,16'd7338,16'd140,16'd6386,16'd1640,16'd6577,16'd1906,-16'd7465,16'd4845,-16'd4988,16'd813,-16'd4065,16'd1064,-16'd7439,16'd2980,16'd468,16'd876,-16'd2020,-16'd6504,-16'd5861,-16'd2140,16'd538,-16'd5514,-16'd6091,16'd2175,-16'd6542,16'd6113,-16'd2741,16'd3216,16'd6508,16'd1341};
dout[383]={ 16'd5123,16'd368,16'd5137,16'd9394,-16'd9444,-16'd11949,-16'd4335,16'd5701,-16'd1759,-16'd2276,16'd4927,16'd1151,-16'd6699,16'd6492,-16'd5428,16'd5418,16'd4015,16'd7157,16'd407,-16'd5537,-16'd1950,-16'd4270,16'd4472,-16'd839,-16'd8753,16'd6101,16'd6714,16'd1780,-16'd2429,-16'd5389,-16'd6674,-16'd3167,-16'd6244,16'd4753,-16'd600,-16'd5843};
dout[384]={ 16'd5266,-16'd5990,-16'd2018,16'd6951,16'd2115,16'd7471,-16'd5055,16'd365,-16'd2990,-16'd6058,-16'd6384,16'd2459,-16'd1696,-16'd3740,-16'd3862,16'd1257,16'd4901,-16'd2250,-16'd5735,16'd384,-16'd6562,16'd5068,16'd4008,-16'd5162,-16'd7212,16'd7636,-16'd2860,16'd3083,-16'd1246,16'd218,16'd8723,16'd623,16'd4642,-16'd2176,16'd7432,-16'd599};
dout[385]={ -16'd1739,16'd4013,-16'd2512,16'd6935,16'd3889,-16'd3535,16'd4579,-16'd2268,-16'd3329,-16'd219,-16'd202,16'd4074,16'd2333,16'd3091,16'd2310,-16'd4596,16'd592,16'd1234,16'd4070,16'd2891,-16'd5473,16'd855,16'd3501,16'd1746,16'd1832,16'd6727,-16'd2915,16'd1154,16'd3128,-16'd1266,-16'd5654,-16'd7437,16'd6909,16'd1533,-16'd4754,-16'd4694};
dout[386]={ 16'd537,-16'd4119,-16'd6119,-16'd732,16'd7008,16'd695,-16'd1770,16'd2779,-16'd3103,-16'd1243,-16'd49,-16'd954,-16'd3392,-16'd4418,16'd5722,16'd3609,16'd2305,-16'd3918,-16'd1712,-16'd609,-16'd1449,-16'd987,16'd3256,-16'd5645,16'd5327,-16'd3849,16'd5235,-16'd5393,16'd6071,16'd490,-16'd2582,16'd4907,16'd4600,16'd4939,-16'd3877,-16'd499};
dout[387]={ -16'd8068,-16'd1772,16'd6115,16'd164,16'd1443,16'd3368,16'd3453,16'd2094,-16'd5251,-16'd2642,16'd4078,16'd3910,-16'd6930,16'd2467,-16'd3102,-16'd900,16'd6456,-16'd7,-16'd3278,-16'd3235,-16'd2283,-16'd4634,-16'd4755,-16'd746,16'd425,16'd1410,-16'd6676,16'd3266,-16'd2340,-16'd2492,-16'd2556,16'd2431,-16'd3118,16'd4466,-16'd1170,-16'd2726};
dout[388]={ -16'd7593,-16'd1249,16'd5264,-16'd710,16'd416,16'd4524,16'd3710,-16'd402,16'd1776,-16'd1137,-16'd6711,16'd2739,-16'd7185,16'd3547,16'd1140,16'd9450,16'd2213,16'd6757,-16'd395,16'd1562,16'd2712,16'd5105,16'd6211,16'd7291,16'd4662,16'd3820,-16'd4028,16'd677,-16'd1674,16'd4740,-16'd3531,-16'd2811,16'd6311,-16'd2552,-16'd4165,-16'd7111};
dout[389]={ -16'd5063,16'd3334,-16'd3205,-16'd4881,-16'd7256,-16'd8899,16'd4524,-16'd2205,16'd5740,16'd1798,-16'd1244,16'd2691,-16'd3553,-16'd810,16'd1561,-16'd3494,16'd484,16'd4236,16'd3987,-16'd6494,16'd104,16'd4831,16'd4037,-16'd1144,16'd2723,16'd1406,16'd5559,-16'd4914,16'd3337,-16'd4452,-16'd2753,16'd3208,16'd453,16'd7820,-16'd4300,-16'd2539};
dout[390]={ -16'd6124,-16'd16589,-16'd5320,16'd5205,16'd1273,16'd6140,16'd1194,-16'd4570,16'd356,-16'd7014,-16'd2731,16'd91,-16'd9137,-16'd6527,16'd2105,-16'd2907,-16'd4017,16'd1584,-16'd1460,16'd4865,-16'd7424,16'd5359,-16'd3596,16'd687,16'd419,16'd10932,16'd7645,16'd7594,16'd3483,-16'd7036,-16'd5169,-16'd743,16'd4771,-16'd2778,-16'd555,16'd1748};
dout[391]={ -16'd834,-16'd7393,16'd4321,-16'd473,16'd1802,16'd1620,16'd4186,16'd5952,-16'd3954,-16'd6647,-16'd841,-16'd2198,-16'd10103,-16'd3007,-16'd5609,16'd6523,16'd4344,16'd6730,16'd2529,16'd611,-16'd9711,-16'd6495,-16'd2918,-16'd262,-16'd2120,16'd8712,-16'd4749,16'd2558,-16'd2159,16'd9505,-16'd10066,16'd2347,-16'd1441,-16'd6826,-16'd7456,-16'd9023};
dout[392]={ 16'd7047,16'd1547,-16'd3864,-16'd333,-16'd913,-16'd4348,-16'd2123,-16'd2624,16'd5578,16'd1667,16'd8052,-16'd2955,16'd2555,-16'd3005,-16'd11251,16'd159,16'd2390,16'd9828,-16'd5389,-16'd1249,-16'd128,-16'd7025,16'd7023,16'd284,16'd6494,-16'd1376,-16'd3132,-16'd3345,-16'd3870,16'd5487,-16'd10269,-16'd3575,-16'd5736,-16'd7299,16'd4809,-16'd6049};
dout[393]={ 16'd2490,-16'd736,-16'd4331,16'd2376,-16'd9006,-16'd5139,16'd1021,-16'd4840,16'd4836,-16'd142,16'd5002,-16'd2993,-16'd219,16'd4788,16'd548,16'd6420,16'd1114,16'd5052,-16'd866,-16'd1698,16'd2444,-16'd8246,-16'd4703,-16'd3821,16'd3723,16'd8683,16'd7967,-16'd6624,-16'd717,-16'd2885,-16'd2966,16'd4550,-16'd2641,-16'd7287,-16'd1307,-16'd3854};
dout[394]={ -16'd3515,-16'd4060,16'd3349,16'd12003,16'd2262,16'd5183,-16'd7073,16'd3575,16'd3272,16'd6588,-16'd5142,16'd155,16'd1357,-16'd5357,-16'd6152,16'd7516,-16'd5849,16'd4699,16'd6736,-16'd2447,-16'd6293,16'd2941,-16'd766,-16'd2171,16'd3771,-16'd446,-16'd6587,-16'd2013,16'd4199,16'd3919,16'd1394,-16'd2950,-16'd3715,-16'd7161,16'd4236,-16'd1247};
dout[395]={ 16'd5503,-16'd9918,-16'd7576,16'd932,-16'd3498,16'd5059,16'd7098,16'd5816,-16'd5850,16'd6237,16'd1613,16'd4899,-16'd4181,16'd2156,-16'd5529,16'd4621,16'd5415,-16'd7099,16'd2258,16'd5911,16'd3796,16'd2077,-16'd8125,-16'd3478,-16'd4302,16'd6891,-16'd5230,16'd1567,16'd3929,-16'd3632,-16'd6366,16'd2347,-16'd2365,-16'd3931,-16'd2090,-16'd2339};
dout[396]={ -16'd8038,-16'd4888,-16'd2898,16'd6497,16'd4507,-16'd1300,16'd5196,16'd665,-16'd3685,16'd7006,-16'd4595,-16'd3322,-16'd660,16'd2851,16'd2528,16'd3151,16'd892,-16'd1005,16'd2988,16'd874,-16'd1019,-16'd2484,-16'd8337,-16'd827,16'd7181,16'd6177,-16'd4210,16'd1876,-16'd7240,16'd6518,-16'd6507,-16'd6183,16'd4485,-16'd6794,-16'd6655,16'd623};
dout[397]={ -16'd4167,-16'd6888,16'd2691,16'd4016,-16'd3807,16'd4489,16'd3538,-16'd4007,-16'd17,-16'd2719,16'd2087,16'd6431,-16'd5932,-16'd7137,-16'd2207,16'd4155,-16'd5195,16'd5864,16'd1795,-16'd5493,-16'd689,16'd5409,-16'd3566,16'd2823,-16'd1762,-16'd1781,16'd1123,16'd4049,-16'd6128,16'd137,-16'd6805,-16'd444,16'd944,16'd601,16'd2871,-16'd6916};
dout[398]={ -16'd4258,-16'd6899,-16'd2976,-16'd2510,16'd5016,16'd900,16'd7353,16'd1159,16'd2248,-16'd356,16'd7935,16'd3409,-16'd9093,-16'd5786,16'd3663,-16'd3449,-16'd1995,-16'd3567,-16'd6154,-16'd367,-16'd3720,-16'd1780,16'd795,16'd521,-16'd4303,-16'd4298,16'd4862,16'd2318,-16'd6742,16'd2435,16'd3589,-16'd34,16'd6615,-16'd1958,16'd4028,16'd3791};
dout[399]={ 16'd1685,16'd5733,16'd51,16'd5221,-16'd1348,-16'd7314,16'd1932,16'd682,16'd266,16'd23,-16'd5113,16'd5674,-16'd859,-16'd3123,-16'd3011,16'd8790,16'd4163,16'd2629,-16'd7393,-16'd6926,16'd7627,-16'd5631,-16'd436,-16'd4407,-16'd598,16'd1823,-16'd845,16'd6306,16'd4459,16'd6776,-16'd2635,16'd671,16'd1291,-16'd2919,-16'd1548,-16'd5630};
dout[400]={ 16'd2875,-16'd16515,-16'd602,-16'd2373,-16'd5728,-16'd1783,16'd6411,16'd378,-16'd4968,-16'd6704,16'd5736,16'd3148,16'd1464,-16'd8049,16'd7405,-16'd118,-16'd11126,-16'd5389,-16'd2715,16'd6729,16'd3578,16'd5842,-16'd2321,-16'd5571,16'd8527,16'd6917,16'd8140,16'd4461,-16'd7387,16'd5216,-16'd3257,-16'd6856,16'd6616,-16'd518,-16'd4592,-16'd6752};
dout[401]={ 16'd3109,16'd2819,16'd3188,-16'd7089,-16'd1948,16'd3862,16'd4476,-16'd6209,16'd1484,-16'd7743,-16'd1074,16'd2067,-16'd3371,16'd8025,-16'd7570,-16'd884,-16'd5256,-16'd3914,16'd6106,16'd8237,-16'd10414,16'd1857,-16'd1713,16'd3033,16'd2666,16'd10078,-16'd3529,16'd4890,-16'd157,16'd2216,16'd1174,-16'd5852,-16'd3101,-16'd10765,16'd6710,-16'd1422};
dout[402]={ 16'd5028,-16'd3474,16'd5472,16'd4400,-16'd5318,-16'd6194,-16'd8132,16'd8381,-16'd2235,-16'd5153,-16'd1281,16'd393,-16'd445,16'd5975,-16'd2555,-16'd10232,16'd4561,-16'd2609,16'd5613,-16'd5577,-16'd5901,16'd4511,-16'd8016,16'd1151,16'd7789,-16'd2794,-16'd1858,-16'd7482,-16'd10757,16'd5926,-16'd7035,16'd1745,-16'd44,-16'd8794,-16'd19,-16'd3501};
dout[403]={ 16'd598,16'd3463,16'd911,16'd6142,16'd4830,-16'd4553,-16'd3634,16'd5633,16'd6476,-16'd4723,16'd2159,-16'd6129,16'd3954,16'd1276,-16'd5949,-16'd4590,16'd10203,16'd1973,16'd5929,16'd3611,-16'd933,-16'd113,-16'd9065,-16'd121,-16'd2679,16'd9330,16'd10380,16'd191,-16'd5625,-16'd602,16'd4374,-16'd6495,16'd370,-16'd4566,-16'd1481,16'd5529};
dout[404]={ -16'd4545,-16'd8716,-16'd8230,-16'd3297,16'd5570,16'd3071,-16'd7435,16'd3913,-16'd4580,-16'd3087,-16'd8178,-16'd6530,-16'd8527,16'd7750,16'd2772,16'd1867,16'd3175,-16'd2262,16'd1770,-16'd3204,-16'd6404,-16'd769,-16'd5705,16'd3226,-16'd5293,16'd9063,-16'd2399,-16'd8396,-16'd4293,-16'd6008,16'd1376,-16'd373,16'd2526,-16'd8661,-16'd2398,-16'd7165};
dout[405]={ 16'd5881,16'd5055,-16'd6130,16'd1203,-16'd1141,16'd3332,16'd788,-16'd6045,-16'd4606,16'd3466,-16'd3997,-16'd2466,16'd3362,16'd2237,16'd2711,16'd6184,-16'd7245,-16'd2736,-16'd5885,16'd706,-16'd6320,-16'd2776,16'd3126,-16'd2059,16'd2222,16'd5479,-16'd128,16'd2781,-16'd7910,-16'd1144,16'd3301,-16'd4088,16'd6517,16'd4967,-16'd2595,16'd250};
dout[406]={ -16'd404,-16'd3373,16'd4877,-16'd5560,16'd1820,16'd343,-16'd5766,-16'd4080,16'd1595,16'd1715,-16'd5613,-16'd1322,-16'd7770,-16'd2003,-16'd2780,16'd3784,-16'd6040,-16'd6544,-16'd4348,-16'd2776,16'd1176,-16'd2957,16'd2373,-16'd3606,-16'd1060,-16'd6464,16'd3630,16'd4382,-16'd5482,-16'd32,-16'd4410,16'd3525,16'd2125,-16'd2373,-16'd740,-16'd2796};
dout[407]={ 16'd5000,16'd593,16'd5359,16'd2804,-16'd430,-16'd2817,16'd6306,16'd8771,-16'd520,16'd834,16'd976,-16'd336,16'd152,16'd2688,16'd3152,16'd1067,16'd4718,-16'd890,16'd1418,-16'd2950,16'd2784,16'd3882,-16'd6218,-16'd5006,16'd2762,16'd1814,16'd4535,-16'd676,16'd702,-16'd790,-16'd5691,16'd5255,16'd7604,-16'd6093,-16'd900,16'd4059};
dout[408]={ 16'd3634,-16'd6605,16'd1823,-16'd3548,-16'd3781,16'd4213,-16'd4275,16'd7414,16'd3796,-16'd5938,16'd150,16'd1775,-16'd4107,-16'd5450,16'd1083,16'd1016,16'd4486,16'd3994,16'd4794,-16'd6384,16'd4421,16'd2170,16'd5093,16'd3727,-16'd505,16'd3182,-16'd2055,-16'd2939,16'd2425,-16'd7113,-16'd1350,16'd4038,-16'd3222,-16'd9519,-16'd1040,-16'd6363};
dout[409]={ -16'd1202,16'd1210,-16'd8256,-16'd3961,16'd3440,-16'd1472,-16'd7027,-16'd5402,16'd6920,-16'd2906,-16'd3520,16'd2542,-16'd771,-16'd7420,-16'd3212,-16'd875,16'd3740,16'd7500,16'd3140,-16'd2521,16'd702,-16'd1101,-16'd5941,-16'd2598,16'd3614,16'd6040,-16'd8438,-16'd5572,-16'd4349,16'd2916,-16'd311,16'd5676,16'd6211,-16'd5641,16'd7539,-16'd2492};
dout[410]={ -16'd4052,-16'd14650,-16'd2761,16'd1567,-16'd317,16'd7818,-16'd9624,16'd8370,-16'd5532,-16'd1872,-16'd598,16'd7907,-16'd4220,-16'd527,16'd10290,16'd5876,-16'd3235,-16'd9980,16'd5685,16'd5319,16'd8187,-16'd6029,16'd699,16'd5745,16'd1740,-16'd6757,16'd6532,-16'd2887,-16'd8376,16'd2492,16'd128,-16'd3281,16'd12228,-16'd1584,16'd6436,16'd41};
dout[411]={ 16'd5589,16'd7780,16'd5446,-16'd2256,16'd4913,-16'd1769,-16'd5365,-16'd1805,-16'd2615,16'd4594,16'd4206,16'd2690,-16'd9398,-16'd2686,16'd4021,-16'd3390,16'd282,16'd5848,-16'd3639,16'd2035,16'd690,16'd1950,-16'd7018,16'd63,16'd8765,16'd4139,16'd6697,16'd3672,-16'd10293,-16'd2511,16'd4040,-16'd6868,16'd3740,16'd589,-16'd4282,-16'd9485};
dout[412]={ -16'd5699,16'd8165,-16'd2393,16'd6127,-16'd10047,-16'd9109,16'd3874,16'd1470,16'd2849,-16'd8343,16'd5425,16'd2175,-16'd7522,16'd823,-16'd6656,-16'd12687,16'd789,-16'd4534,16'd4861,16'd4998,-16'd9415,16'd1237,16'd6419,-16'd5648,16'd2215,-16'd5276,-16'd3993,-16'd4358,-16'd3342,16'd7267,-16'd3832,-16'd4734,16'd5905,-16'd5409,16'd4266,-16'd4350};
dout[413]={ 16'd4290,-16'd5201,16'd5467,-16'd2836,16'd4027,-16'd6332,-16'd1431,-16'd1379,-16'd5582,16'd6331,16'd290,16'd2278,-16'd8820,-16'd4388,16'd4304,-16'd6089,16'd3107,16'd1827,-16'd8490,16'd1268,-16'd4911,-16'd576,16'd2887,-16'd8344,16'd241,-16'd3861,16'd5599,-16'd9039,16'd5711,-16'd2861,16'd302,-16'd4661,-16'd35,16'd3323,-16'd5030,16'd5525};
dout[414]={ -16'd271,-16'd2211,-16'd6381,16'd5316,16'd4809,16'd5208,-16'd4330,-16'd6135,16'd5217,-16'd2225,-16'd1188,-16'd5875,16'd965,16'd5139,-16'd2261,16'd7851,-16'd4380,16'd2564,-16'd8628,16'd4578,-16'd6575,16'd3783,-16'd8368,-16'd2073,-16'd7734,16'd1714,16'd8512,16'd1941,-16'd1866,-16'd3366,-16'd6719,-16'd1879,-16'd5235,16'd4218,16'd628,16'd4534};
dout[415]={ -16'd782,-16'd6583,-16'd4447,16'd1571,-16'd3395,16'd2772,-16'd7941,-16'd8709,-16'd7087,16'd6155,16'd3698,-16'd3245,16'd1696,-16'd564,16'd8219,-16'd650,-16'd5650,16'd2279,-16'd672,16'd5789,16'd152,-16'd8140,-16'd8170,-16'd1289,-16'd386,-16'd2269,-16'd1223,-16'd6618,-16'd1764,16'd4213,-16'd3,-16'd5631,-16'd2348,-16'd2284,16'd901,16'd1717};
dout[416]={ 16'd2377,16'd5242,16'd2988,-16'd2503,16'd4018,-16'd5127,16'd1335,16'd4014,16'd238,16'd973,-16'd3694,16'd566,-16'd5165,16'd127,16'd2966,16'd5706,-16'd1431,-16'd3308,16'd1307,-16'd5224,16'd1803,16'd3282,16'd367,16'd5177,-16'd1948,-16'd6571,-16'd3795,16'd2800,-16'd1469,-16'd5034,-16'd5115,16'd2421,16'd620,16'd5504,-16'd3557,16'd4948};
dout[417]={ 16'd2859,-16'd2076,-16'd2389,16'd5117,16'd6911,16'd5843,-16'd7151,16'd2844,-16'd5172,16'd4510,16'd2423,16'd2353,16'd5805,-16'd4003,-16'd1720,16'd4453,-16'd2081,16'd8113,16'd289,16'd626,-16'd1508,16'd5229,16'd40,-16'd5074,-16'd1622,16'd2780,-16'd124,-16'd1605,16'd6497,16'd5985,16'd7125,16'd5807,16'd794,-16'd4965,16'd3482,16'd4910};
dout[418]={ -16'd4056,-16'd2911,16'd4334,-16'd6747,-16'd5153,16'd968,-16'd6219,-16'd3631,16'd2243,16'd8055,16'd9216,16'd619,16'd5574,-16'd3873,16'd5749,-16'd2224,-16'd1674,-16'd840,16'd4639,16'd114,16'd5522,16'd4977,16'd3068,16'd904,-16'd6519,-16'd5984,16'd3326,-16'd6764,16'd4997,16'd1833,16'd1484,16'd2616,-16'd1605,16'd1357,-16'd4842,16'd2210};
dout[419]={ -16'd3168,-16'd2842,-16'd7125,-16'd1943,16'd3696,-16'd7738,-16'd7944,-16'd6132,16'd3856,16'd3336,16'd8208,16'd284,16'd1410,-16'd6219,16'd328,16'd3757,16'd2022,-16'd1112,-16'd3868,-16'd2488,16'd2029,-16'd2003,-16'd4097,-16'd7955,-16'd8661,16'd5196,-16'd5190,-16'd682,16'd2515,-16'd4878,-16'd4901,16'd5710,-16'd743,-16'd1530,-16'd2963,-16'd994};
dout[420]={ 16'd5426,16'd685,16'd2826,16'd4374,16'd4439,16'd2987,-16'd9546,16'd4867,-16'd3237,16'd3077,-16'd742,16'd2061,-16'd8784,-16'd2971,16'd6494,16'd10584,-16'd9302,-16'd871,-16'd1858,16'd6500,16'd1607,16'd1860,-16'd2994,-16'd8474,16'd9022,-16'd8347,16'd9480,-16'd8736,-16'd7545,16'd3446,-16'd3265,16'd498,16'd8272,-16'd6195,16'd1255,-16'd1248};
dout[421]={ -16'd4982,16'd10515,16'd6616,16'd3959,16'd7178,16'd5084,-16'd1519,-16'd7227,16'd5111,-16'd8604,-16'd857,16'd1335,16'd3569,16'd8721,16'd560,-16'd9261,-16'd4719,-16'd781,16'd5136,16'd8687,16'd1295,-16'd5858,-16'd3939,-16'd3139,16'd696,16'd6302,16'd1963,-16'd3249,-16'd5769,16'd5862,-16'd1927,-16'd4584,16'd9339,-16'd3070,16'd4220,-16'd5971};
dout[422]={ -16'd8201,16'd6058,-16'd2247,16'd5445,-16'd7304,-16'd3311,-16'd6724,16'd2449,16'd7652,16'd2860,-16'd3258,16'd3421,-16'd9638,16'd4155,-16'd223,-16'd7127,-16'd7887,16'd6950,-16'd8237,-16'd2632,-16'd4156,-16'd5234,-16'd3390,16'd3854,16'd6439,16'd1160,16'd4758,-16'd7062,-16'd8519,16'd5408,-16'd3151,-16'd8633,16'd7899,-16'd8411,16'd6553,-16'd2103};
dout[423]={ -16'd6213,-16'd3798,16'd1843,16'd5674,16'd389,-16'd7673,16'd2202,-16'd6317,16'd7044,-16'd2290,-16'd349,-16'd6506,-16'd7734,-16'd6373,16'd7291,16'd529,-16'd1724,16'd4160,-16'd2949,-16'd611,-16'd5512,-16'd9235,-16'd1575,-16'd3958,16'd992,16'd5261,16'd13182,-16'd7444,-16'd2971,16'd1422,16'd8619,-16'd10689,16'd2244,16'd1409,-16'd3645,-16'd3244};
dout[424]={ 16'd2147,-16'd4672,16'd4320,16'd5718,-16'd2628,-16'd3099,-16'd1587,16'd2931,16'd5685,-16'd5606,-16'd2459,-16'd182,16'd5620,-16'd2297,16'd10285,-16'd4174,16'd9180,-16'd1440,-16'd6044,-16'd2605,16'd4790,16'd5867,-16'd9671,16'd2221,-16'd579,-16'd6064,-16'd473,-16'd10845,16'd1220,-16'd6477,-16'd6351,-16'd7606,16'd3141,16'd2275,-16'd2321,-16'd1596};
dout[425]={ -16'd6948,-16'd2719,16'd1465,-16'd5866,16'd4376,16'd3977,16'd5907,-16'd3735,-16'd1472,-16'd2547,-16'd5629,-16'd3625,16'd6950,16'd5890,16'd4995,16'd252,-16'd2097,16'd2270,-16'd1450,-16'd3487,16'd7669,16'd3279,-16'd7580,-16'd2304,-16'd6838,-16'd9282,16'd5340,-16'd5533,16'd4962,-16'd271,16'd7644,16'd5009,-16'd1742,-16'd2711,16'd391,-16'd7253};
dout[426]={ 16'd2887,16'd1271,-16'd3764,-16'd2568,-16'd7667,16'd2065,-16'd1783,16'd5552,-16'd4403,16'd770,16'd2765,-16'd1809,16'd3338,-16'd2113,-16'd4807,-16'd3554,16'd3272,16'd4090,-16'd4051,-16'd3023,16'd6247,-16'd3302,16'd226,-16'd5598,16'd4110,-16'd3404,-16'd892,-16'd6879,-16'd7417,16'd885,-16'd554,16'd2013,16'd6642,-16'd4757,-16'd4013,16'd5747};
dout[427]={ -16'd795,16'd3685,-16'd6543,-16'd2544,16'd5299,-16'd165,-16'd4430,16'd4204,16'd2708,-16'd3009,-16'd5191,16'd2964,16'd6615,-16'd7344,-16'd711,16'd7364,-16'd4560,-16'd1160,16'd1966,-16'd265,-16'd1913,-16'd1256,16'd1612,-16'd1936,16'd3896,-16'd3334,-16'd4709,-16'd2081,-16'd2109,16'd5751,-16'd2383,-16'd2554,-16'd746,16'd718,16'd374,-16'd445};
dout[428]={ 16'd6430,16'd1094,16'd2253,16'd4192,16'd1231,-16'd884,-16'd309,-16'd5108,-16'd1222,-16'd590,16'd4876,16'd1685,-16'd8190,-16'd10112,16'd4511,-16'd689,16'd3770,16'd111,16'd3624,-16'd8153,-16'd1215,-16'd1303,-16'd4044,16'd5485,-16'd368,16'd6781,16'd1774,-16'd982,-16'd1014,-16'd305,16'd1074,16'd7976,-16'd6501,16'd3199,16'd5335,-16'd3768};
dout[429]={ 16'd1058,-16'd3423,-16'd238,16'd4045,-16'd65,16'd159,16'd1555,-16'd4771,-16'd3388,16'd1051,16'd1383,-16'd2484,-16'd2873,-16'd6534,-16'd6129,16'd4164,-16'd4313,-16'd1913,-16'd3168,-16'd7474,-16'd5665,-16'd869,16'd2104,-16'd2879,-16'd2653,-16'd362,16'd1030,16'd789,16'd7256,16'd3958,16'd9034,16'd3963,-16'd611,-16'd5427,16'd6086,16'd2032};
dout[430]={ 16'd1969,-16'd4010,16'd6886,16'd269,16'd2250,16'd4840,16'd4705,16'd6741,-16'd5002,-16'd190,16'd6029,-16'd214,-16'd4511,-16'd1952,-16'd51,-16'd29,-16'd12733,-16'd3165,16'd1425,16'd970,16'd2602,-16'd6007,16'd2938,-16'd1118,16'd7349,-16'd18740,-16'd1853,-16'd5580,-16'd502,16'd792,16'd7634,16'd7172,16'd3951,-16'd4785,16'd2674,-16'd4056};
dout[431]={ 16'd7020,16'd4861,-16'd3478,-16'd5494,16'd3329,16'd933,16'd1474,-16'd2000,-16'd416,-16'd684,16'd3298,16'd850,-16'd6233,16'd5364,-16'd575,-16'd2737,16'd1916,16'd4679,-16'd5747,-16'd4540,16'd6332,-16'd9033,-16'd1447,16'd1904,16'd5520,-16'd4435,16'd8086,-16'd6391,-16'd4515,-16'd332,-16'd7651,-16'd7879,16'd4020,-16'd1615,-16'd4033,-16'd6};
dout[432]={ -16'd660,16'd5008,-16'd3954,16'd2430,-16'd8759,-16'd1089,16'd5876,16'd4743,16'd1889,-16'd3271,-16'd4898,-16'd5243,-16'd3743,16'd411,16'd1752,-16'd14379,16'd1812,16'd5538,16'd419,16'd6773,-16'd1428,16'd2505,-16'd2329,-16'd1673,16'd5638,16'd7095,-16'd2973,-16'd8728,-16'd7264,16'd9302,-16'd9214,-16'd5609,16'd8435,-16'd7314,16'd6293,-16'd2731};
dout[433]={ -16'd236,16'd1302,-16'd62,-16'd749,16'd3657,16'd5054,16'd3764,-16'd7384,16'd4008,-16'd2586,16'd4410,16'd6078,-16'd5602,-16'd1070,16'd6875,-16'd9142,-16'd4219,-16'd5252,16'd622,-16'd5264,16'd6388,-16'd6624,16'd7065,-16'd8883,16'd2281,-16'd5591,16'd9417,-16'd8766,-16'd4652,-16'd5322,-16'd543,-16'd7849,-16'd4125,16'd743,-16'd4037,16'd53};
dout[434]={ 16'd6113,-16'd4458,16'd6825,-16'd6814,16'd7059,16'd1435,-16'd5358,-16'd5546,16'd6887,-16'd3144,-16'd1180,16'd2115,-16'd7667,16'd5031,16'd4027,16'd5478,16'd3270,16'd251,-16'd7201,-16'd6407,16'd4801,16'd3263,-16'd5467,16'd4825,16'd2186,-16'd270,16'd4067,-16'd4789,-16'd1838,-16'd5200,-16'd6176,16'd1918,-16'd311,16'd6339,16'd2869,-16'd785};
dout[435]={ -16'd3599,-16'd1111,-16'd4234,-16'd7721,16'd1489,-16'd3829,-16'd4730,-16'd5867,-16'd8973,-16'd2920,16'd642,-16'd6072,-16'd8671,16'd5316,16'd4691,16'd3995,16'd5369,-16'd1270,-16'd5549,-16'd3296,-16'd497,-16'd5871,16'd3645,-16'd6653,-16'd4726,-16'd10538,16'd1577,16'd732,-16'd3198,16'd950,-16'd2804,16'd5371,-16'd4069,-16'd3583,-16'd2363,-16'd4039};
dout[436]={ 16'd5522,-16'd2601,16'd118,16'd4052,16'd4572,16'd2695,-16'd6765,16'd5304,-16'd234,-16'd2523,-16'd4848,16'd5383,-16'd3240,-16'd5206,16'd1005,16'd35,16'd2739,16'd2958,-16'd3158,16'd1367,-16'd3145,-16'd4003,-16'd3805,-16'd7013,-16'd2528,16'd7044,-16'd4856,-16'd8612,16'd5621,16'd1319,-16'd1733,16'd4008,16'd2966,16'd2051,16'd4763,16'd4815};
dout[437]={ 16'd3310,16'd5722,16'd7002,16'd2071,-16'd287,-16'd6128,16'd2321,-16'd872,-16'd179,-16'd5466,16'd5493,-16'd930,-16'd503,-16'd6152,16'd2952,-16'd486,-16'd1724,16'd3810,16'd128,16'd3121,16'd5761,16'd526,-16'd4257,16'd2840,-16'd1388,-16'd5992,-16'd4965,16'd924,-16'd3008,-16'd6176,-16'd1429,16'd4527,-16'd4961,-16'd1251,-16'd397,16'd859};
dout[438]={ 16'd4044,-16'd4187,-16'd5861,-16'd3959,-16'd1743,16'd4051,16'd2876,16'd817,16'd5862,-16'd2809,-16'd4474,16'd41,16'd2073,16'd1478,-16'd7521,16'd6297,-16'd5323,16'd7914,16'd764,-16'd4178,16'd4858,-16'd453,16'd321,16'd492,-16'd5763,16'd5121,16'd5686,-16'd4709,-16'd2115,-16'd5563,16'd2202,16'd2268,16'd219,-16'd112,16'd4503,16'd7176};
dout[439]={ 16'd868,16'd7682,-16'd5854,16'd7007,-16'd1177,-16'd2574,-16'd430,-16'd1449,-16'd1937,16'd918,16'd6444,-16'd714,-16'd6944,-16'd6129,16'd3968,-16'd2023,16'd6795,16'd777,-16'd2600,16'd2816,-16'd507,16'd5053,16'd734,16'd2473,-16'd5963,16'd2972,-16'd7197,-16'd115,16'd5104,16'd5645,-16'd3132,-16'd1057,-16'd2137,16'd10151,-16'd227,-16'd3706};
dout[440]={ -16'd5585,-16'd1207,16'd1861,16'd1018,-16'd3357,16'd5858,-16'd3041,-16'd5849,16'd2079,16'd1908,16'd2403,16'd9353,-16'd7698,-16'd554,-16'd4121,-16'd2651,-16'd6956,-16'd12848,16'd285,-16'd8627,16'd2861,16'd2239,-16'd7043,-16'd7388,16'd8596,-16'd6778,-16'd8661,-16'd2577,16'd6707,-16'd7244,-16'd2889,16'd95,16'd13403,16'd3067,-16'd2188,16'd7345};
dout[441]={ 16'd899,16'd10105,16'd534,16'd9646,16'd985,16'd8061,16'd8413,16'd2684,-16'd3509,-16'd3898,-16'd3547,-16'd6522,-16'd5399,-16'd2250,16'd3556,-16'd7250,16'd512,-16'd176,-16'd2284,16'd6094,16'd8708,-16'd8270,16'd4268,16'd3042,-16'd3142,16'd4791,16'd1014,-16'd1475,-16'd1453,-16'd1542,16'd5121,-16'd5674,-16'd2438,-16'd1273,16'd309,-16'd3043};
dout[442]={ -16'd3735,16'd6120,-16'd7277,-16'd3146,-16'd2214,16'd5716,16'd36,-16'd7524,16'd4027,-16'd3147,16'd2558,16'd4597,16'd1916,-16'd1537,-16'd914,-16'd10850,16'd1854,16'd3426,-16'd4802,-16'd4416,16'd3121,16'd404,16'd7250,16'd442,16'd6041,16'd7924,16'd2753,-16'd33,-16'd6514,16'd5220,-16'd539,16'd924,16'd1354,-16'd2068,16'd3125,-16'd4093};
dout[443]={ -16'd3204,-16'd2050,-16'd1200,-16'd4263,-16'd1265,16'd4233,16'd1305,16'd519,16'd3935,-16'd7780,-16'd4941,16'd524,16'd1074,-16'd11841,16'd2717,16'd4343,16'd2917,-16'd2091,16'd6028,16'd1297,16'd9984,16'd1241,16'd3060,-16'd4884,16'd6699,-16'd4397,16'd4265,16'd413,16'd1677,16'd7104,16'd6642,16'd6043,-16'd1843,-16'd4738,-16'd8751,16'd8310};
dout[444]={ 16'd6625,16'd3410,-16'd3253,-16'd1990,-16'd1997,-16'd7766,16'd5042,16'd272,16'd6528,-16'd1982,-16'd1755,16'd5759,-16'd5326,-16'd2338,-16'd3589,16'd1487,16'd6617,16'd3288,16'd2415,16'd2157,16'd8295,16'd664,-16'd5818,-16'd2683,-16'd3462,-16'd4381,16'd7182,-16'd1112,16'd1205,-16'd5567,-16'd3977,16'd2404,16'd250,-16'd333,16'd8142,16'd1229};
dout[445]={ -16'd5256,16'd3588,16'd4198,-16'd1245,-16'd7740,16'd5897,-16'd1893,16'd2538,16'd2153,16'd3329,-16'd1072,16'd4309,-16'd6064,16'd3324,-16'd7855,-16'd4332,-16'd7005,16'd2689,-16'd7740,-16'd2260,-16'd1236,-16'd6811,16'd985,-16'd4398,16'd3758,-16'd5289,16'd1989,-16'd8687,16'd4544,-16'd4768,16'd2514,16'd7494,-16'd7220,-16'd810,16'd5561,16'd6538};
dout[446]={ 16'd6398,-16'd5196,-16'd6631,-16'd4338,-16'd6388,16'd3549,-16'd6076,16'd3670,16'd271,-16'd4613,-16'd1444,-16'd2291,16'd1365,16'd5631,-16'd5651,-16'd414,-16'd5242,-16'd78,-16'd6647,-16'd247,-16'd7277,16'd18,16'd8696,16'd1899,16'd3172,-16'd3510,16'd6958,16'd3536,16'd2013,-16'd2830,16'd7932,16'd3337,-16'd2759,16'd584,16'd2786,-16'd2158};
dout[447]={ 16'd7651,16'd1311,-16'd125,-16'd5260,-16'd1508,16'd2498,16'd4096,-16'd2583,-16'd3592,16'd533,16'd5384,16'd1983,-16'd7563,-16'd369,-16'd6200,-16'd4016,-16'd2991,-16'd2740,-16'd2820,-16'd1961,-16'd5220,-16'd6999,-16'd2502,-16'd5104,16'd1101,16'd7325,16'd1493,16'd4933,-16'd1509,16'd5108,16'd6595,16'd4516,16'd500,16'd7219,16'd1574,16'd787};
dout[448]={ 16'd3943,16'd8750,16'd668,-16'd2156,-16'd977,16'd5666,16'd4580,-16'd6688,16'd7823,-16'd5816,-16'd1166,16'd1128,-16'd7410,16'd2290,-16'd7140,16'd298,-16'd5105,-16'd4769,16'd3403,-16'd79,16'd4079,-16'd2467,-16'd2065,-16'd1018,-16'd1966,16'd644,16'd795,-16'd5292,-16'd4049,16'd362,-16'd4578,-16'd5897,-16'd767,16'd8539,-16'd2672,-16'd1055};
dout[449]={ 16'd2959,16'd1298,16'd3103,16'd6051,16'd5376,-16'd6455,16'd1989,-16'd6963,16'd3130,16'd1219,16'd3089,-16'd4958,16'd2293,-16'd7897,-16'd473,16'd2408,16'd5972,16'd5658,16'd4451,-16'd627,-16'd5977,-16'd2341,-16'd3943,-16'd7994,16'd1514,16'd5259,-16'd1680,-16'd6744,16'd4215,16'd5107,16'd3969,16'd4560,-16'd4303,-16'd1007,-16'd6981,16'd5626};
dout[450]={ 16'd710,-16'd1593,16'd1647,16'd9911,-16'd6996,16'd5457,16'd6785,16'd744,16'd11579,-16'd1519,16'd1390,16'd2441,16'd2104,16'd399,-16'd1142,-16'd1782,-16'd7755,-16'd7031,-16'd6170,-16'd9346,-16'd9899,-16'd5001,16'd9884,16'd3788,-16'd1863,-16'd10005,-16'd7558,-16'd8550,-16'd4149,-16'd10465,16'd6676,16'd2173,16'd4955,16'd6353,16'd831,-16'd6205};
dout[451]={ -16'd4909,16'd5508,16'd2721,16'd4206,-16'd2391,16'd947,16'd4730,16'd199,16'd735,-16'd2907,-16'd2026,16'd2798,-16'd9997,16'd4957,-16'd3511,-16'd1013,16'd4297,-16'd1858,-16'd6731,-16'd1500,16'd2306,-16'd4508,16'd5443,-16'd1137,-16'd3356,-16'd3370,16'd971,16'd872,-16'd1660,16'd2383,-16'd4558,-16'd1130,16'd6948,-16'd7629,-16'd3037,-16'd1376};
dout[452]={ 16'd4963,16'd1929,-16'd4689,-16'd4455,-16'd7822,16'd7664,-16'd636,16'd622,16'd1634,16'd2652,-16'd3632,-16'd3993,-16'd9473,-16'd4199,-16'd5422,-16'd5860,16'd4264,-16'd3610,-16'd3297,16'd4677,16'd5611,-16'd9307,16'd6437,16'd2776,16'd2697,16'd2236,-16'd6240,-16'd6983,-16'd7041,16'd8443,-16'd5626,-16'd766,-16'd1012,-16'd3505,-16'd461,-16'd2386};
dout[453]={ 16'd9216,16'd5924,16'd3768,16'd3805,-16'd9685,-16'd154,-16'd5027,-16'd8800,16'd4020,-16'd6349,-16'd1364,16'd1203,16'd4015,-16'd4101,-16'd2537,-16'd7486,16'd6152,-16'd5733,-16'd4925,16'd498,16'd5455,16'd4274,-16'd4962,16'd1590,16'd1737,16'd849,-16'd1119,-16'd6656,16'd4125,16'd4126,16'd1410,16'd2849,-16'd9660,-16'd2437,16'd2902,-16'd2250};
dout[454]={ 16'd3405,16'd2925,-16'd1848,16'd6692,-16'd5083,16'd502,-16'd2483,-16'd1666,-16'd611,16'd5107,16'd8377,-16'd1287,-16'd6481,16'd4729,-16'd8806,-16'd5537,16'd2215,-16'd2669,-16'd6392,-16'd1743,16'd2150,-16'd5584,-16'd2314,16'd1594,16'd10385,-16'd2575,16'd5593,-16'd4580,16'd456,16'd2280,16'd5029,16'd1282,-16'd11055,-16'd1740,16'd1953,16'd5435};
dout[455]={ -16'd723,16'd4622,-16'd1898,-16'd522,-16'd1446,-16'd5711,16'd7639,-16'd6246,-16'd5889,-16'd186,-16'd1403,16'd1452,-16'd1748,16'd4093,-16'd10835,-16'd1443,-16'd2756,-16'd7245,16'd5658,16'd4262,16'd3973,-16'd2113,16'd5865,-16'd619,-16'd2906,-16'd2722,16'd6193,16'd238,-16'd5427,16'd2050,-16'd993,-16'd2937,-16'd2409,-16'd258,16'd6595,16'd1660};
dout[456]={ 16'd2946,16'd3715,-16'd7791,16'd858,16'd1144,16'd3567,-16'd3648,16'd3155,16'd22,-16'd6340,16'd6288,16'd6502,-16'd1547,-16'd2596,-16'd3488,16'd9187,16'd6562,-16'd7367,16'd479,16'd2899,16'd4218,16'd198,16'd167,16'd2517,-16'd5606,-16'd4215,-16'd862,16'd4575,16'd1307,16'd1635,16'd1381,-16'd1499,-16'd5732,-16'd2874,-16'd71,-16'd1184};
dout[457]={ 16'd2389,16'd2457,-16'd1737,-16'd5052,-16'd1992,16'd4757,16'd5063,16'd3185,-16'd2263,16'd7926,-16'd1524,16'd4975,-16'd3224,16'd4894,16'd2823,-16'd3513,-16'd3510,16'd5314,16'd4184,16'd4880,-16'd576,-16'd6873,-16'd3510,-16'd6195,-16'd3087,16'd4783,-16'd4207,-16'd1492,16'd7075,-16'd2779,-16'd5962,-16'd2320,16'd2713,-16'd5173,-16'd1246,-16'd5452};
dout[458]={ -16'd4234,-16'd1465,16'd3429,16'd2398,16'd6971,16'd2446,-16'd4170,-16'd3198,16'd1413,-16'd6037,16'd2057,-16'd2838,-16'd617,-16'd6918,-16'd3916,-16'd7157,16'd6350,16'd4189,-16'd4333,16'd5981,16'd1101,-16'd4490,16'd3640,16'd2062,-16'd6886,16'd1927,-16'd674,-16'd5426,16'd4161,16'd1361,16'd3694,-16'd5073,-16'd6308,-16'd2317,-16'd5741,16'd2477};
dout[459]={ 16'd7544,16'd744,16'd8117,16'd6773,16'd1944,16'd2773,-16'd4368,16'd838,16'd860,-16'd2683,-16'd4200,-16'd3094,16'd5261,-16'd8397,16'd1305,-16'd1499,16'd2139,16'd2495,-16'd7999,-16'd2654,16'd6089,16'd6193,16'd3496,-16'd6444,-16'd14,16'd6036,-16'd34,-16'd5768,16'd3364,-16'd2113,-16'd5687,16'd4210,16'd4290,16'd4610,16'd4178,16'd5296};
dout[460]={ 16'd794,16'd4915,-16'd5608,16'd829,16'd1674,16'd2803,-16'd3322,16'd6252,16'd11847,-16'd7617,16'd3868,16'd2162,-16'd6662,-16'd5673,-16'd7195,16'd6133,-16'd2477,16'd2702,16'd500,-16'd11762,-16'd7996,16'd4739,16'd9193,-16'd7581,16'd5584,-16'd10348,-16'd3690,-16'd2247,-16'd2080,-16'd7243,-16'd2291,-16'd5648,16'd3385,16'd3843,16'd2542,16'd5405};
dout[461]={ 16'd5408,16'd6494,16'd3279,-16'd4350,-16'd11324,16'd116,16'd7247,-16'd3528,-16'd3881,-16'd2430,16'd805,-16'd7657,-16'd4542,16'd5776,16'd5681,-16'd8815,-16'd6961,-16'd2820,-16'd4517,-16'd5009,16'd9199,-16'd9160,-16'd1028,-16'd6357,-16'd3628,16'd7182,-16'd6182,-16'd4059,16'd2349,16'd292,16'd2215,16'd943,16'd7570,-16'd3182,-16'd4813,-16'd7530};
dout[462]={ 16'd7514,16'd6649,16'd1518,-16'd206,-16'd1814,16'd144,16'd1637,16'd2996,-16'd9261,16'd1986,-16'd1795,16'd1760,-16'd5258,16'd10528,-16'd2896,-16'd4496,-16'd176,16'd2031,16'd2285,-16'd7021,-16'd1136,-16'd1056,-16'd1732,16'd3968,16'd4205,-16'd3536,-16'd15356,16'd252,-16'd10498,16'd2243,-16'd964,16'd9120,16'd6928,16'd1037,-16'd5326,-16'd2421};
dout[463]={ 16'd1459,-16'd4069,16'd4113,-16'd4193,-16'd2129,-16'd7825,16'd5921,16'd2708,16'd587,-16'd2824,16'd8763,16'd8142,-16'd3547,-16'd5648,16'd5833,16'd4661,16'd6927,-16'd1492,16'd632,-16'd6690,-16'd2964,16'd4380,16'd1000,16'd3339,16'd2035,-16'd7354,16'd105,-16'd2524,-16'd4872,16'd1786,16'd870,16'd2121,-16'd3642,-16'd3054,16'd4102,-16'd3879};
dout[464]={ 16'd8403,-16'd6859,-16'd5547,16'd4315,16'd674,-16'd6804,16'd390,-16'd2326,16'd6600,-16'd4235,16'd8599,16'd3400,-16'd8215,-16'd7366,16'd4750,16'd1414,-16'd4137,-16'd6425,16'd2301,16'd4770,16'd1135,16'd5560,16'd7760,16'd2084,16'd696,16'd5496,16'd1089,16'd954,16'd448,-16'd4520,-16'd2567,16'd5203,-16'd9959,-16'd504,-16'd1054,16'd1418};
dout[465]={ -16'd7198,16'd1029,-16'd8594,-16'd4811,-16'd3837,16'd787,16'd2561,-16'd1779,16'd1800,-16'd3822,16'd7792,16'd4525,-16'd8587,16'd1390,-16'd1459,-16'd2253,16'd2439,16'd6560,-16'd5307,-16'd3800,-16'd3874,-16'd7561,-16'd3424,16'd2279,16'd7222,-16'd7731,-16'd5595,16'd4335,16'd5901,-16'd1098,-16'd4111,16'd5139,-16'd2411,-16'd5490,-16'd6829,16'd1242};
dout[466]={ 16'd3526,16'd1082,-16'd8138,-16'd792,-16'd7386,16'd3198,16'd2162,-16'd356,16'd3986,16'd1423,-16'd5769,16'd5594,-16'd5602,16'd1707,16'd3363,-16'd4178,16'd1830,16'd6416,-16'd6865,16'd4548,-16'd6379,-16'd7155,-16'd4425,-16'd4336,16'd6692,16'd8656,-16'd2824,-16'd4493,16'd2624,16'd3576,-16'd3293,-16'd3447,16'd3683,16'd2753,16'd7854,16'd2045};
dout[467]={ -16'd2726,-16'd1222,16'd4300,16'd7298,-16'd3039,-16'd4101,-16'd4857,16'd2726,-16'd5316,-16'd2477,16'd3001,-16'd7495,-16'd2177,16'd3686,16'd3122,-16'd3575,16'd2967,16'd3838,-16'd2179,-16'd1113,-16'd3821,-16'd1525,16'd6609,16'd47,16'd3249,-16'd3275,16'd7291,-16'd481,16'd6845,-16'd4060,-16'd783,16'd5185,16'd780,-16'd3741,-16'd2762,-16'd1699};
dout[468]={ -16'd576,-16'd844,-16'd1389,-16'd6621,16'd6607,16'd646,-16'd2458,-16'd3989,16'd834,-16'd1107,-16'd5056,-16'd5082,-16'd4632,-16'd8501,-16'd836,-16'd978,-16'd2326,-16'd5331,16'd2672,-16'd4428,16'd4382,16'd2161,16'd750,16'd1009,-16'd3933,-16'd3201,16'd882,16'd3255,16'd3595,-16'd2945,16'd7552,-16'd3112,-16'd4090,-16'd2661,-16'd1934,16'd3528};
dout[469]={ -16'd227,16'd7094,-16'd2487,-16'd5900,-16'd4031,16'd1118,16'd227,-16'd412,16'd5952,16'd6576,-16'd210,-16'd1238,-16'd4440,-16'd3573,16'd7457,-16'd6259,16'd4039,-16'd4416,-16'd4563,16'd6463,-16'd7144,16'd4163,-16'd4505,-16'd3498,16'd3877,16'd2876,16'd3457,16'd2414,16'd5644,-16'd4815,-16'd1062,-16'd8843,16'd4188,-16'd7660,16'd3869,16'd1547};
dout[470]={ -16'd4266,-16'd6268,-16'd909,16'd7401,-16'd8755,-16'd7920,-16'd4512,-16'd1186,-16'd792,-16'd1124,16'd7224,16'd4077,16'd3345,16'd2496,16'd2328,16'd4860,-16'd6109,16'd18,16'd4299,-16'd10513,-16'd9455,16'd1124,16'd4045,16'd2384,-16'd4845,-16'd9211,-16'd395,16'd6203,-16'd922,-16'd10323,16'd1190,-16'd3497,16'd2858,16'd5192,16'd6112,-16'd8538};
dout[471]={ 16'd217,16'd595,-16'd8544,-16'd6829,-16'd1340,16'd312,-16'd2637,16'd7353,16'd4180,-16'd9685,-16'd1681,-16'd1799,16'd4547,16'd3094,16'd724,-16'd7169,-16'd2391,-16'd2902,16'd2006,-16'd8809,-16'd2247,-16'd8395,16'd602,-16'd2138,16'd5465,16'd7607,-16'd12107,-16'd2114,-16'd6453,-16'd1032,-16'd1420,16'd5523,16'd5279,16'd5795,-16'd6044,-16'd5794};
dout[472]={ 16'd4609,-16'd1961,16'd2626,16'd4768,-16'd10387,16'd1512,-16'd4660,-16'd9239,-16'd7558,-16'd6288,-16'd175,16'd3774,16'd223,-16'd1232,16'd5250,-16'd7035,-16'd5615,16'd6951,16'd5041,-16'd2267,16'd4362,-16'd8489,16'd5363,-16'd78,-16'd5937,16'd1223,-16'd2135,-16'd934,-16'd8892,16'd7897,-16'd6701,16'd4900,16'd7352,-16'd2280,16'd4093,-16'd2995};
dout[473]={ -16'd743,16'd7278,16'd74,-16'd1010,-16'd9434,-16'd2202,16'd897,-16'd3350,-16'd3979,16'd3129,16'd6957,16'd5505,-16'd1161,16'd2406,16'd6699,-16'd2678,-16'd1522,16'd9735,-16'd4936,16'd3748,16'd1034,-16'd6807,16'd1755,-16'd5271,16'd2172,-16'd6219,-16'd558,-16'd6478,16'd1579,-16'd4755,-16'd4979,-16'd1024,-16'd2616,16'd55,-16'd280,16'd2162};
dout[474]={ 16'd7023,16'd2889,16'd4635,16'd3496,16'd3209,-16'd8451,-16'd3916,16'd3028,16'd9348,16'd5437,16'd5400,16'd256,16'd6634,-16'd3762,16'd4696,16'd9613,-16'd2188,16'd6704,16'd2094,-16'd4390,-16'd1279,-16'd7408,-16'd2846,16'd1078,-16'd747,-16'd2814,16'd2686,16'd6145,-16'd4936,-16'd863,-16'd5107,16'd274,-16'd463,16'd2990,16'd2123,16'd766};
dout[475]={ -16'd2746,16'd533,-16'd8857,-16'd4672,16'd493,-16'd7729,-16'd1891,-16'd7624,-16'd1006,16'd172,16'd131,16'd2220,16'd1893,16'd1968,-16'd1298,16'd1211,-16'd1793,-16'd4028,-16'd7024,-16'd3923,16'd3199,-16'd924,16'd4207,16'd4441,16'd6582,16'd669,16'd6942,-16'd3456,16'd2985,-16'd1245,-16'd6749,-16'd4149,-16'd3467,-16'd5606,-16'd2993,16'd6673};
dout[476]={ 16'd3890,16'd3202,16'd3739,16'd5958,-16'd7781,-16'd5830,-16'd5483,16'd273,-16'd1235,-16'd636,16'd3520,16'd2553,16'd3660,-16'd3340,-16'd675,-16'd2882,16'd4799,-16'd2449,16'd4858,-16'd1940,-16'd7126,16'd7786,-16'd643,-16'd4991,16'd245,16'd2639,16'd2265,16'd5307,-16'd4599,16'd1190,-16'd5012,16'd1747,-16'd3214,16'd2670,-16'd2839,-16'd5318};
dout[477]={ -16'd674,16'd5758,-16'd12118,16'd2962,16'd5395,-16'd3650,-16'd5730,16'd3520,-16'd611,16'd384,16'd4722,16'd4026,16'd3529,16'd4485,-16'd2843,16'd6317,-16'd994,-16'd3418,-16'd3776,16'd204,-16'd3363,-16'd4788,16'd350,16'd462,-16'd4713,16'd8718,-16'd712,16'd4855,-16'd5756,-16'd5068,-16'd4457,-16'd877,16'd3707,16'd8362,-16'd1469,16'd1718};
dout[478]={ 16'd1249,16'd4826,-16'd6445,-16'd7797,16'd2702,-16'd2820,-16'd943,-16'd5747,-16'd7180,16'd5283,16'd2586,-16'd6663,-16'd6571,16'd4202,16'd5482,-16'd3910,-16'd2179,16'd6806,-16'd7374,16'd6239,-16'd5707,-16'd4029,-16'd2555,16'd2261,16'd4711,-16'd283,-16'd5146,16'd3087,-16'd3407,-16'd7284,16'd7114,-16'd3066,-16'd6443,-16'd5655,-16'd4844,16'd2467};
dout[479]={ 16'd7078,-16'd2479,-16'd8303,16'd3034,-16'd5062,16'd10068,-16'd3609,-16'd1863,16'd2338,16'd930,-16'd504,16'd5189,16'd1400,-16'd6442,-16'd1900,-16'd6770,-16'd5092,16'd4380,-16'd1968,16'd1589,-16'd94,16'd151,16'd1712,-16'd8082,-16'd1719,16'd3333,16'd1224,-16'd7723,-16'd7993,-16'd2403,16'd1984,16'd1439,16'd5568,16'd2147,-16'd4424,-16'd708};
dout[480]={ -16'd5954,16'd110,16'd3163,16'd7855,-16'd5414,-16'd8383,16'd2593,-16'd4345,16'd7675,-16'd774,16'd3404,16'd8143,-16'd3353,16'd5448,-16'd2716,16'd1191,16'd773,16'd4087,-16'd2060,-16'd11551,-16'd1592,-16'd9224,-16'd9465,-16'd1870,-16'd6691,16'd6470,-16'd8571,-16'd1430,-16'd4196,-16'd9340,-16'd3009,-16'd6058,16'd4778,16'd4744,16'd8973,-16'd7452};
dout[481]={ -16'd4902,16'd4729,16'd1092,-16'd4846,-16'd6492,-16'd2011,-16'd2693,16'd1188,-16'd749,16'd1771,16'd6824,16'd2714,16'd1403,16'd3188,16'd457,-16'd1180,-16'd4165,-16'd1004,-16'd6692,-16'd1357,16'd1222,16'd3297,-16'd1127,-16'd4854,-16'd3961,-16'd1998,-16'd8712,16'd5560,-16'd1249,16'd8940,-16'd2486,-16'd2551,16'd343,-16'd4021,-16'd7612,-16'd5533};
dout[482]={ 16'd7461,16'd7294,16'd6648,-16'd2885,-16'd9405,16'd6453,16'd666,-16'd2895,-16'd12501,-16'd5004,16'd7394,16'd4227,-16'd1532,16'd5344,-16'd7237,-16'd6059,16'd1902,-16'd1701,-16'd930,-16'd8977,16'd6036,16'd5191,16'd5258,-16'd1692,16'd202,16'd5321,16'd1308,-16'd6681,-16'd4566,-16'd286,-16'd5348,-16'd1687,16'd3918,16'd342,16'd3053,16'd4794};
dout[483]={ 16'd7968,-16'd3554,16'd1549,-16'd5184,-16'd449,-16'd6280,16'd2917,-16'd4137,-16'd4698,-16'd3122,16'd6816,16'd10865,16'd283,16'd2520,16'd6726,-16'd2360,16'd6517,16'd11575,-16'd1364,16'd2091,-16'd6290,-16'd7092,-16'd7795,16'd2618,16'd6068,-16'd3370,-16'd11103,-16'd1196,16'd1891,-16'd8360,16'd1910,-16'd6110,16'd8563,-16'd1471,16'd6611,-16'd2476};
dout[484]={ 16'd550,16'd3162,16'd2158,16'd6550,-16'd8982,-16'd2176,-16'd4337,-16'd5371,16'd1888,16'd4720,16'd3571,-16'd3195,-16'd695,-16'd4225,-16'd1488,16'd140,-16'd2359,16'd1738,16'd2757,-16'd2715,-16'd6948,16'd684,16'd2851,-16'd742,-16'd1527,-16'd2949,-16'd6454,16'd2629,16'd6018,-16'd395,16'd2016,16'd3827,16'd361,-16'd6134,16'd9875,16'd4475};
dout[485]={ -16'd5673,-16'd2321,-16'd6440,16'd5659,16'd3411,-16'd5741,-16'd9107,-16'd5312,16'd9251,-16'd7808,16'd5961,16'd5,16'd7190,16'd4643,-16'd4760,16'd4012,16'd2943,16'd2386,-16'd8488,-16'd1471,-16'd5347,16'd3567,-16'd3528,-16'd6928,16'd3843,-16'd4410,-16'd5836,16'd238,16'd686,-16'd1510,-16'd5352,-16'd4854,-16'd1942,-16'd4574,16'd2942,16'd4647};
dout[486]={ -16'd5748,16'd6224,-16'd2026,16'd1760,-16'd4011,-16'd6107,-16'd5142,-16'd4919,-16'd3251,16'd4325,16'd78,16'd5124,-16'd1107,16'd3301,16'd7356,-16'd4526,-16'd7163,16'd1165,16'd887,16'd6357,-16'd2862,16'd6704,16'd1491,-16'd3020,16'd3333,16'd2005,16'd7406,16'd2606,-16'd3241,16'd3821,-16'd2416,16'd1483,-16'd1480,-16'd5783,16'd4027,16'd724};
dout[487]={ 16'd3129,-16'd3428,-16'd1499,-16'd2243,16'd1290,-16'd1525,16'd5976,16'd408,16'd3730,-16'd5844,-16'd1391,-16'd4259,-16'd785,16'd989,-16'd334,16'd3723,-16'd4628,-16'd728,16'd6766,16'd1515,-16'd7110,-16'd4387,-16'd697,-16'd9,16'd4918,-16'd4266,16'd8741,16'd928,-16'd6761,-16'd1768,16'd6381,16'd4059,-16'd3157,-16'd5907,16'd2488,-16'd2103};
dout[488]={ 16'd4653,-16'd3179,-16'd8657,-16'd7801,16'd8002,16'd4106,16'd1798,16'd5144,16'd683,16'd9654,16'd3471,-16'd6015,-16'd6945,16'd1426,-16'd206,16'd691,16'd2426,-16'd1515,16'd5076,16'd7911,-16'd5795,16'd5948,-16'd1649,16'd5973,-16'd765,-16'd578,16'd816,-16'd2066,-16'd3591,-16'd631,16'd3202,16'd3418,16'd3135,-16'd2635,-16'd1048,16'd4976};
dout[489]={ 16'd6264,16'd5200,-16'd6450,16'd1002,16'd2447,16'd3179,16'd1464,-16'd2925,16'd5799,16'd762,-16'd8405,-16'd1391,-16'd2851,16'd5589,-16'd1207,16'd2462,-16'd1538,-16'd4981,16'd3392,16'd5274,-16'd4874,16'd487,16'd4492,-16'd8217,16'd6485,-16'd6121,-16'd757,-16'd2624,16'd361,-16'd2494,16'd5537,-16'd1254,-16'd4057,16'd3082,16'd1870,-16'd1600};
dout[490]={ 16'd2167,16'd5834,16'd7813,16'd7354,-16'd10978,16'd2514,16'd5524,-16'd6454,-16'd5290,-16'd5918,16'd9218,16'd2207,-16'd3509,-16'd191,-16'd6397,16'd1061,-16'd5028,-16'd321,16'd1692,-16'd6077,16'd380,-16'd4213,-16'd13871,16'd220,-16'd1152,-16'd1707,-16'd3357,-16'd4942,-16'd2121,-16'd7216,-16'd7081,-16'd1671,16'd7503,16'd1348,16'd9137,-16'd4448};
dout[491]={ 16'd4401,-16'd1443,16'd3373,-16'd9691,-16'd3243,16'd5033,16'd5989,16'd6748,-16'd4548,16'd172,-16'd2063,-16'd57,-16'd7085,16'd7175,16'd6334,-16'd7886,-16'd1117,16'd5621,-16'd3753,-16'd483,16'd3855,16'd596,-16'd7078,-16'd7437,-16'd2848,16'd1026,-16'd7094,-16'd350,-16'd2970,16'd7780,-16'd2894,-16'd2259,-16'd2537,16'd545,16'd3173,16'd2923};
dout[492]={ -16'd3675,16'd6773,-16'd478,-16'd11948,-16'd12132,16'd277,-16'd1389,16'd5235,-16'd6458,-16'd7167,16'd1478,16'd902,-16'd8322,16'd8356,16'd2190,-16'd916,16'd1408,16'd8874,16'd1615,-16'd2457,16'd1451,-16'd4874,16'd443,16'd3413,16'd3916,-16'd1265,16'd1717,16'd4885,16'd1645,16'd2383,-16'd9800,-16'd3090,16'd542,16'd6274,-16'd473,16'd963};
dout[493]={ 16'd4359,-16'd4225,16'd9282,-16'd2547,-16'd4646,-16'd2054,-16'd693,-16'd3742,-16'd8968,-16'd7090,-16'd896,16'd3308,16'd3819,16'd960,-16'd1191,-16'd428,-16'd3429,16'd8164,16'd5521,16'd3904,-16'd3002,-16'd7088,16'd2476,-16'd63,-16'd5526,-16'd4051,-16'd6294,16'd3128,16'd5994,-16'd2284,16'd301,16'd2099,16'd7052,-16'd680,16'd5280,16'd82};
dout[494]={ -16'd1362,16'd703,-16'd3809,16'd2334,16'd1720,-16'd8122,16'd890,-16'd6715,-16'd2998,16'd6817,-16'd6100,16'd6251,16'd5037,16'd901,-16'd3025,-16'd2417,16'd4268,16'd3355,-16'd7876,-16'd7679,-16'd3953,16'd6421,16'd5078,-16'd6805,16'd5063,-16'd948,-16'd3555,16'd1629,16'd5594,-16'd2064,16'd107,-16'd3845,-16'd1532,16'd4408,16'd8650,-16'd3126};
dout[495]={ -16'd586,-16'd1855,-16'd4185,-16'd4093,16'd481,16'd74,-16'd9106,-16'd1246,16'd2235,-16'd3035,16'd1881,-16'd7687,-16'd7372,-16'd4894,-16'd4920,-16'd31,-16'd1405,16'd6874,16'd3861,16'd1193,-16'd6193,16'd469,-16'd4985,-16'd3243,-16'd5932,-16'd3997,-16'd1211,-16'd4981,-16'd3897,16'd156,16'd1871,16'd7940,16'd3951,16'd600,16'd2833,16'd3295};
dout[496]={ -16'd1251,-16'd4585,-16'd6805,16'd1984,-16'd4022,16'd4606,-16'd5869,16'd1510,16'd7455,16'd247,16'd3890,16'd251,-16'd1509,16'd6683,-16'd3888,16'd4280,16'd3532,-16'd1623,16'd2318,-16'd3464,-16'd7184,16'd3258,-16'd4700,-16'd4455,16'd7607,16'd5128,16'd7414,16'd2741,16'd5479,-16'd661,16'd3289,16'd7322,-16'd5311,16'd1049,-16'd3025,16'd2860};
dout[497]={ -16'd5235,16'd5558,-16'd1147,-16'd5446,16'd2027,16'd1359,16'd3727,-16'd5541,16'd446,-16'd3562,-16'd2343,-16'd6787,-16'd3000,16'd3735,16'd5596,16'd784,-16'd4624,16'd4050,-16'd5082,16'd2251,-16'd5762,16'd402,16'd4848,-16'd3812,-16'd5109,16'd4400,16'd4099,-16'd842,-16'd2610,-16'd3613,16'd7136,16'd4589,16'd2882,-16'd6684,16'd5786,-16'd6480};
dout[498]={ -16'd1999,16'd7154,-16'd7811,-16'd436,-16'd147,16'd6554,16'd2390,16'd2638,16'd2239,16'd8865,-16'd668,16'd3974,-16'd173,16'd1507,16'd2105,16'd4278,-16'd3362,16'd5524,16'd5525,-16'd1855,16'd3278,16'd3412,16'd861,16'd3507,16'd1814,16'd3463,-16'd3219,16'd1331,16'd439,-16'd7902,-16'd6031,-16'd5342,-16'd6515,16'd4325,16'd4214,-16'd6153};
dout[499]={ -16'd1170,-16'd5107,-16'd4380,-16'd261,-16'd3484,-16'd4694,-16'd7280,-16'd7516,-16'd6549,16'd3777,16'd1273,16'd2168,-16'd4343,-16'd5005,-16'd6103,-16'd1197,-16'd5122,-16'd7438,-16'd5361,-16'd1639,16'd4682,-16'd2219,16'd3881,16'd1519,16'd6610,16'd2547,-16'd753,-16'd4836,-16'd5550,-16'd4698,16'd3412,-16'd2802,-16'd4660,-16'd774,-16'd4053,16'd6294};
dout[500]={ 16'd5598,16'd7773,-16'd73,-16'd545,-16'd8300,16'd2060,-16'd5968,-16'd5941,16'd1844,-16'd11828,-16'd489,16'd2791,-16'd5274,-16'd1041,16'd1990,16'd7093,-16'd7410,16'd4715,-16'd4183,-16'd6206,-16'd1072,-16'd6942,-16'd17602,-16'd1527,16'd1748,16'd5411,-16'd7412,-16'd3172,16'd6733,-16'd4687,-16'd1460,-16'd3873,-16'd2667,-16'd2850,16'd1972,16'd5321};
dout[501]={ 16'd2751,-16'd4444,-16'd2081,-16'd5351,-16'd6435,16'd5413,-16'd6258,-16'd1548,-16'd4410,-16'd6784,16'd8398,-16'd5743,-16'd6991,16'd7382,-16'd3683,-16'd5754,-16'd1815,-16'd2058,-16'd4457,-16'd7084,-16'd7785,-16'd7466,-16'd5168,-16'd3614,-16'd1901,-16'd560,16'd1086,-16'd7067,16'd526,16'd1963,16'd1553,16'd802,16'd3499,16'd1593,-16'd4960,-16'd8434};
dout[502]={ -16'd2903,-16'd2549,16'd4921,-16'd11799,-16'd3813,16'd8248,-16'd712,-16'd2381,-16'd37,-16'd7715,16'd7923,16'd4979,-16'd3052,16'd4058,-16'd4505,16'd5410,16'd3323,16'd6297,16'd1397,-16'd1136,-16'd1713,-16'd5879,-16'd1359,-16'd7335,16'd4130,16'd4714,-16'd9622,-16'd5565,16'd6722,-16'd2264,-16'd4923,-16'd6840,-16'd3709,-16'd3020,16'd3284,-16'd2457};
dout[503]={ 16'd5005,-16'd439,16'd6124,-16'd5395,-16'd359,-16'd5526,-16'd3274,16'd5386,-16'd1654,16'd1182,16'd821,16'd6499,16'd3477,16'd7232,16'd3834,16'd4847,16'd6682,16'd5948,-16'd3542,16'd5637,16'd1102,16'd3048,-16'd2606,-16'd8381,-16'd3522,-16'd799,-16'd6210,-16'd145,-16'd2746,-16'd10958,16'd1367,-16'd2719,16'd2455,-16'd2741,16'd8851,-16'd8478};
dout[504]={ -16'd5851,-16'd7970,-16'd259,-16'd4680,-16'd1675,-16'd4651,16'd5913,-16'd4950,16'd2505,16'd3314,-16'd6700,16'd9233,-16'd7869,16'd4005,-16'd2919,-16'd5045,16'd3220,16'd5312,16'd4246,-16'd1162,16'd2278,16'd3659,16'd2919,16'd2743,-16'd5188,16'd3456,-16'd3398,16'd5663,16'd1130,-16'd9332,16'd3136,16'd3766,16'd3067,-16'd8120,16'd6973,16'd5540};
dout[505]={ -16'd5108,16'd1679,16'd361,16'd3916,16'd1347,-16'd686,-16'd7443,16'd2419,-16'd6368,-16'd2904,-16'd2180,16'd5302,-16'd4789,16'd7173,-16'd544,16'd1585,16'd265,-16'd2050,16'd5389,-16'd3181,16'd1218,16'd1839,-16'd4731,-16'd5675,16'd2717,16'd5182,-16'd157,16'd4084,-16'd15,16'd6046,-16'd2993,16'd9442,-16'd3251,16'd4874,16'd3498,16'd1755};
dout[506]={ -16'd642,16'd8412,-16'd1091,-16'd3316,16'd2855,-16'd4837,16'd170,-16'd7282,-16'd4898,-16'd1040,-16'd6108,-16'd3594,-16'd449,-16'd4272,16'd5213,16'd763,-16'd2710,16'd989,16'd4597,16'd6185,16'd2088,16'd591,-16'd1071,-16'd1920,-16'd4798,16'd874,-16'd970,-16'd309,-16'd2711,-16'd2792,16'd723,16'd3270,16'd199,16'd713,-16'd3985,-16'd1769};
dout[507]={ 16'd5072,-16'd1446,16'd5962,16'd4383,-16'd6489,-16'd2252,16'd4013,-16'd8249,-16'd4948,16'd5621,-16'd3608,16'd1792,16'd1544,16'd4571,-16'd2297,16'd2544,-16'd5228,-16'd653,16'd1755,-16'd833,16'd4019,16'd6718,-16'd5785,16'd2329,16'd8396,16'd4445,16'd3728,-16'd4148,-16'd2398,-16'd4999,16'd778,16'd1691,16'd3668,-16'd2823,16'd4940,16'd1613};
dout[508]={ -16'd1635,-16'd4515,-16'd6052,-16'd2449,-16'd93,16'd4193,-16'd8604,16'd24,-16'd574,-16'd413,16'd2786,-16'd6465,16'd1046,16'd7468,16'd2600,-16'd7646,16'd880,16'd3494,-16'd220,-16'd5487,16'd5897,-16'd2591,16'd4027,-16'd5047,-16'd2918,-16'd2458,16'd7232,16'd7315,16'd7374,16'd5265,16'd2938,16'd6358,16'd371,16'd1561,16'd263,-16'd7343};
dout[509]={ -16'd217,-16'd4792,-16'd2544,-16'd24,16'd4324,16'd8427,16'd3365,-16'd3753,-16'd5088,-16'd4299,16'd1737,-16'd3600,16'd6012,16'd1121,16'd1791,16'd3737,16'd3519,16'd7955,16'd5222,16'd359,-16'd4345,-16'd2669,16'd6205,-16'd3258,16'd4332,-16'd5313,16'd605,-16'd6774,16'd1443,-16'd4219,16'd3010,16'd3775,-16'd5197,16'd6461,16'd3949,-16'd5928};
dout[510]={ -16'd295,-16'd1418,-16'd40,16'd2595,-16'd4829,-16'd3813,16'd4010,-16'd4882,16'd5479,-16'd8812,-16'd1316,16'd5810,16'd1864,-16'd4354,16'd1467,16'd7287,-16'd219,-16'd6712,16'd4450,16'd11304,16'd1933,-16'd6430,-16'd11819,-16'd2810,16'd3616,-16'd6235,16'd243,16'd6219,-16'd2100,-16'd371,-16'd2577,16'd7180,-16'd2678,16'd3824,16'd9597,16'd5779};
dout[511]={ 16'd3172,16'd3251,-16'd1120,16'd2803,16'd376,-16'd1646,16'd171,-16'd4208,16'd900,16'd4709,-16'd3790,-16'd4979,16'd5131,-16'd4161,-16'd7776,-16'd3279,-16'd8062,16'd2461,-16'd4779,-16'd3740,16'd4899,16'd4116,-16'd439,-16'd9451,16'd1889,-16'd852,-16'd5042,-16'd1094,-16'd1938,-16'd24,16'd2940,16'd295,-16'd1134,16'd8351,-16'd229,16'd5386};
dout[512]={ 16'd6365,16'd3179,-16'd5038,-16'd4690,-16'd4284,16'd2079,-16'd613,16'd1426,16'd855,-16'd5110,16'd2567,-16'd9208,16'd3957,16'd1504,-16'd6056,16'd2307,16'd1159,16'd9516,-16'd2794,16'd4167,-16'd5644,-16'd5060,16'd5661,-16'd9607,-16'd2835,16'd1869,-16'd9800,-16'd817,16'd1239,16'd9150,16'd2226,16'd21,-16'd5036,-16'd849,16'd2445,-16'd6845};
dout[513]={ 16'd5163,-16'd403,-16'd1284,-16'd10023,16'd2133,-16'd1211,16'd8745,16'd4301,16'd3114,16'd7674,-16'd9877,16'd1291,16'd869,-16'd1129,16'd4638,16'd7065,-16'd3943,-16'd2123,-16'd4436,-16'd5604,-16'd5810,-16'd6584,-16'd7095,16'd2830,16'd2012,16'd230,-16'd1866,16'd2712,16'd8047,-16'd1712,-16'd7119,-16'd3744,16'd3638,16'd3940,16'd1260,16'd5101};
dout[514]={ 16'd4918,-16'd3671,16'd10120,16'd201,-16'd6928,-16'd1484,-16'd4934,-16'd3420,16'd3744,16'd10856,-16'd14220,16'd4946,-16'd6761,16'd3570,16'd6134,-16'd5686,-16'd3329,16'd1145,16'd1878,16'd2192,16'd91,-16'd6522,16'd6777,-16'd4260,-16'd5852,-16'd4981,16'd3776,16'd1823,16'd1322,-16'd800,-16'd1268,16'd3530,-16'd6309,16'd792,16'd1356,-16'd8107};
dout[515]={ 16'd1823,16'd7120,16'd6819,16'd1752,-16'd7596,16'd4783,-16'd6863,-16'd6618,-16'd857,16'd2223,16'd3254,-16'd2436,16'd4487,-16'd4972,-16'd1484,16'd58,-16'd6634,-16'd3356,-16'd1416,16'd3892,-16'd4501,-16'd2338,16'd5885,16'd4729,-16'd2133,16'd7933,16'd5189,16'd4401,16'd4118,-16'd1321,-16'd3490,16'd9652,16'd4006,-16'd7501,16'd3307,-16'd2360};
dout[516]={ -16'd1878,-16'd1510,-16'd3595,16'd379,16'd4684,16'd6382,-16'd7280,-16'd3077,-16'd3060,-16'd5742,16'd4690,16'd3928,-16'd3811,16'd4758,-16'd5537,16'd6055,-16'd3225,16'd9893,-16'd5984,-16'd6536,16'd4537,16'd1172,16'd8111,16'd4127,16'd8307,-16'd2455,16'd963,16'd5899,-16'd6695,-16'd236,16'd2642,-16'd3276,16'd4807,-16'd1588,16'd5306,16'd4414};
dout[517]={ 16'd536,-16'd1989,16'd272,16'd2953,-16'd4904,16'd3419,-16'd6278,-16'd6242,16'd407,-16'd2002,-16'd7160,16'd1646,-16'd4534,-16'd4194,-16'd5673,-16'd2909,16'd125,-16'd5403,-16'd6801,-16'd571,-16'd2406,16'd4865,16'd3959,-16'd8197,16'd5155,-16'd1174,16'd1019,16'd6073,16'd2691,16'd2264,16'd2325,-16'd911,-16'd1773,16'd2593,16'd3584,-16'd2573};
dout[518]={ -16'd2368,-16'd5106,-16'd1026,16'd2084,-16'd1570,-16'd990,-16'd1109,-16'd4430,16'd407,-16'd5710,-16'd1039,-16'd7738,-16'd752,-16'd2361,16'd5810,16'd1807,-16'd5423,16'd5528,16'd3698,-16'd1172,-16'd2410,16'd4629,-16'd5187,16'd2314,-16'd4590,16'd980,16'd412,-16'd1697,-16'd5366,-16'd5499,-16'd5427,16'd674,16'd6996,-16'd4515,16'd2716,-16'd6523};
dout[519]={ -16'd4598,-16'd1122,-16'd1358,16'd1228,-16'd1302,-16'd4555,-16'd3330,-16'd4942,-16'd6167,16'd1053,-16'd7643,-16'd988,16'd4496,16'd6115,16'd4251,16'd4883,16'd3888,-16'd1800,16'd2680,16'd7262,16'd4063,16'd3213,16'd3699,16'd1872,-16'd1463,-16'd3801,-16'd5861,-16'd2,-16'd1781,-16'd444,16'd277,16'd3634,16'd5061,-16'd6997,16'd276,16'd5859};
dout[520]={ 16'd5950,16'd1674,-16'd2578,16'd6134,-16'd2997,-16'd1517,16'd6501,-16'd5056,-16'd5618,16'd3012,-16'd1343,16'd11828,16'd4320,-16'd31,-16'd6482,16'd11128,-16'd4332,-16'd8287,16'd5356,16'd1939,-16'd2786,-16'd4556,-16'd13587,16'd1489,16'd9781,16'd3214,-16'd3572,16'd7147,-16'd404,-16'd6307,-16'd433,-16'd5165,-16'd8852,16'd7235,16'd8715,16'd6357};
dout[521]={ 16'd1223,16'd3477,-16'd1604,16'd1775,-16'd2607,16'd1786,16'd7305,-16'd7631,16'd965,16'd1318,-16'd280,-16'd3284,-16'd4030,16'd791,16'd3848,-16'd6822,16'd2191,16'd8728,-16'd3852,16'd3889,-16'd1432,-16'd427,-16'd993,16'd1145,16'd6107,-16'd3218,-16'd6835,-16'd1079,-16'd4584,16'd8994,-16'd5615,-16'd1810,16'd110,16'd6398,16'd3464,-16'd1250};
dout[522]={ -16'd2054,16'd7893,16'd3907,-16'd5341,-16'd5174,-16'd5074,-16'd4084,-16'd7768,-16'd2278,16'd4021,16'd6007,-16'd11825,16'd5783,-16'd6042,-16'd8751,16'd3286,-16'd2066,16'd5842,-16'd6493,-16'd1675,-16'd5453,-16'd4790,-16'd969,16'd2976,-16'd7251,-16'd1834,-16'd5577,16'd450,16'd156,16'd4041,-16'd4819,-16'd7723,-16'd2385,16'd3275,-16'd3985,-16'd4347};
dout[523]={ 16'd6370,16'd1600,16'd4751,-16'd8886,-16'd6285,-16'd7154,16'd4440,16'd2034,-16'd1257,-16'd1714,16'd332,-16'd4015,16'd2798,16'd5691,-16'd3041,-16'd3735,-16'd4444,16'd1464,-16'd8434,16'd1505,-16'd1992,-16'd148,-16'd5630,-16'd2641,-16'd1472,16'd1438,16'd5850,16'd8438,-16'd5180,-16'd7018,-16'd4628,-16'd194,-16'd8738,16'd4368,16'd8410,16'd3908};
dout[524]={ 16'd1068,-16'd5667,16'd6071,16'd4631,-16'd7365,-16'd6447,16'd2104,16'd6611,16'd3325,-16'd622,-16'd7928,16'd1383,16'd1862,16'd8921,-16'd3473,16'd1156,16'd1633,16'd817,-16'd3308,16'd6237,-16'd8222,-16'd8206,16'd680,16'd1822,-16'd4559,16'd3671,16'd1531,16'd421,-16'd2644,16'd498,-16'd6098,16'd8282,-16'd7843,-16'd3530,-16'd2176,16'd3200};
dout[525]={ -16'd4905,-16'd7946,16'd9061,-16'd10277,-16'd6203,-16'd4431,-16'd5560,16'd3204,-16'd7013,16'd949,-16'd5440,16'd5850,-16'd3207,16'd2814,-16'd2629,-16'd3021,16'd2312,16'd665,16'd4542,16'd6674,-16'd1489,-16'd7271,-16'd107,16'd2379,-16'd1185,-16'd6131,-16'd2186,16'd5016,16'd5155,-16'd2090,-16'd6826,-16'd1930,16'd596,-16'd1332,-16'd6405,-16'd4048};
dout[526]={ -16'd1381,16'd7187,16'd7458,16'd1925,-16'd585,-16'd1666,-16'd6215,16'd288,-16'd730,16'd6209,-16'd1264,16'd3383,-16'd2706,-16'd4443,-16'd969,16'd254,16'd2296,16'd4889,-16'd5707,-16'd4913,16'd3227,-16'd6259,16'd7627,-16'd367,-16'd122,-16'd7019,-16'd577,16'd6356,-16'd5341,16'd1655,16'd212,-16'd141,-16'd1542,-16'd6784,-16'd7509,-16'd815};
dout[527]={ 16'd3812,16'd1847,16'd5345,-16'd5114,-16'd4525,16'd3697,-16'd8010,-16'd6790,16'd3750,16'd7266,16'd4400,-16'd1090,-16'd7410,16'd512,16'd2519,16'd5251,-16'd980,-16'd5174,-16'd4316,-16'd3980,-16'd971,-16'd1486,-16'd6032,-16'd3155,16'd682,16'd2871,-16'd1042,-16'd964,-16'd6413,-16'd875,16'd4257,16'd1065,-16'd939,16'd4995,16'd5033,-16'd8792};
dout[528]={ -16'd5968,16'd3009,-16'd2667,-16'd3663,16'd1338,-16'd6106,-16'd3184,-16'd5850,-16'd2467,-16'd5193,-16'd850,16'd4147,16'd5170,16'd5426,16'd5721,-16'd7396,-16'd3150,-16'd460,16'd554,16'd1916,-16'd4400,-16'd2168,-16'd20,-16'd4298,16'd3821,16'd203,16'd2166,-16'd1471,-16'd1451,16'd5236,16'd3593,-16'd2234,16'd1611,-16'd490,16'd2556,-16'd3342};
dout[529]={ 16'd4537,-16'd5000,16'd3759,-16'd558,16'd668,16'd6790,-16'd4056,16'd4803,16'd6707,-16'd4644,-16'd3031,-16'd5415,-16'd1142,16'd3095,-16'd6264,-16'd7734,16'd3849,16'd5258,16'd7178,16'd4099,16'd427,-16'd1915,-16'd499,-16'd219,16'd5031,16'd2430,16'd4988,16'd752,16'd5494,16'd427,16'd3657,16'd5165,16'd2440,16'd5003,16'd164,-16'd2359};
dout[530]={ -16'd251,16'd1236,-16'd2129,-16'd1155,16'd4388,-16'd469,-16'd4201,-16'd5863,16'd186,-16'd1033,-16'd4469,16'd6146,16'd6312,-16'd10655,16'd2211,16'd268,-16'd6423,16'd3899,-16'd7683,-16'd1596,-16'd978,16'd579,-16'd191,-16'd2056,16'd6556,-16'd2099,16'd5590,16'd4773,16'd5686,16'd2460,16'd1139,-16'd1573,16'd3633,16'd6215,-16'd185,16'd1632};
dout[531]={ -16'd29,16'd63,-16'd4138,-16'd6524,-16'd4560,16'd5374,16'd4960,16'd680,-16'd3279,-16'd3460,-16'd7238,-16'd7494,-16'd218,-16'd5431,-16'd5236,-16'd4923,-16'd5340,-16'd1997,16'd4396,16'd7209,-16'd5035,16'd2845,-16'd8001,16'd5709,16'd5841,16'd4117,-16'd6449,-16'd5846,16'd6123,16'd972,-16'd3531,16'd5689,-16'd6071,16'd2428,16'd2318,-16'd2622};
dout[532]={ 16'd8663,16'd370,-16'd10200,16'd2819,16'd1244,16'd7178,-16'd3402,16'd5274,-16'd1010,16'd10025,16'd1312,-16'd1781,-16'd7012,-16'd4896,16'd4471,16'd4767,16'd3328,-16'd3226,-16'd322,16'd2210,-16'd1447,16'd1735,-16'd4820,16'd3993,16'd7769,-16'd8634,-16'd1506,-16'd5207,16'd3287,16'd9258,-16'd9780,16'd3939,-16'd4571,-16'd2125,16'd5630,16'd2553};
dout[533]={ -16'd3586,-16'd2114,-16'd2654,-16'd3992,16'd3354,16'd4655,-16'd5279,16'd3871,-16'd8918,16'd7940,-16'd8319,16'd1052,-16'd7804,-16'd1507,-16'd3041,16'd6738,16'd4792,-16'd7310,-16'd4935,-16'd1436,16'd1345,-16'd7089,-16'd2566,-16'd5523,-16'd404,16'd4382,16'd4734,16'd3090,16'd741,16'd3923,16'd1743,-16'd4129,16'd668,16'd168,-16'd5673,-16'd3809};
dout[534]={ -16'd2532,16'd2968,-16'd2339,-16'd2285,16'd3401,-16'd5263,16'd1649,-16'd2957,16'd6633,-16'd5257,-16'd13245,16'd6712,16'd445,16'd1812,16'd5680,16'd3330,16'd4877,16'd152,16'd2267,16'd514,-16'd393,-16'd690,16'd2013,-16'd1216,-16'd5210,-16'd4557,-16'd2627,16'd822,16'd1144,-16'd7599,-16'd2591,16'd1629,-16'd1079,-16'd1269,-16'd7720,-16'd9480};
dout[535]={ -16'd2452,16'd3115,-16'd479,-16'd3609,16'd2979,16'd184,16'd5662,-16'd4345,16'd6340,16'd2139,-16'd5241,16'd1053,-16'd6307,-16'd4574,16'd6069,16'd2882,-16'd7330,-16'd410,-16'd3626,-16'd1432,16'd3031,-16'd753,-16'd3867,16'd5320,-16'd3410,-16'd6652,16'd869,16'd5087,16'd5551,-16'd4870,16'd3190,-16'd3290,-16'd5212,16'd1020,-16'd2090,-16'd3258};
dout[536]={ -16'd1906,16'd1606,16'd723,16'd705,-16'd7888,-16'd1389,16'd1101,16'd1838,16'd5991,16'd2673,16'd2465,16'd985,-16'd3786,16'd4938,16'd6265,16'd142,-16'd4304,16'd1790,16'd4925,16'd6469,16'd1105,-16'd8294,16'd4086,16'd1788,-16'd4367,16'd4729,-16'd6225,-16'd1094,-16'd2564,-16'd2868,-16'd1726,16'd1039,-16'd4934,16'd4284,-16'd6529,-16'd1168};
dout[537]={ 16'd2841,-16'd1416,16'd514,-16'd5447,-16'd4358,-16'd1920,-16'd2452,-16'd4959,-16'd5040,16'd7181,-16'd3641,-16'd2999,-16'd6855,16'd4629,-16'd5306,16'd2162,-16'd1601,-16'd5844,16'd3704,16'd3631,-16'd2849,16'd1776,16'd2546,-16'd8371,16'd3709,-16'd977,16'd1099,-16'd5153,16'd2553,-16'd4588,16'd695,-16'd3787,-16'd2275,16'd2911,-16'd3362,-16'd7435};
dout[538]={ 16'd5026,-16'd2306,16'd4930,16'd7263,16'd6536,16'd2422,-16'd2247,16'd1788,-16'd394,-16'd78,-16'd1260,-16'd2397,16'd1707,-16'd658,16'd165,-16'd5297,-16'd4129,-16'd7245,-16'd1247,-16'd2528,16'd3999,-16'd6394,16'd3506,-16'd7320,-16'd6081,-16'd4748,16'd143,16'd3506,-16'd1163,-16'd1724,-16'd729,16'd2844,-16'd6487,-16'd230,16'd3525,-16'd2827};
dout[539]={ -16'd1855,16'd1569,16'd1984,-16'd1869,16'd3862,16'd6186,-16'd5548,-16'd4768,16'd5762,16'd4076,-16'd5843,16'd3887,16'd2813,16'd1543,16'd608,16'd5116,16'd1933,-16'd5257,-16'd1300,16'd5565,16'd3053,16'd1979,16'd5390,16'd2539,16'd3327,-16'd1202,16'd6598,-16'd6393,16'd4614,16'd125,-16'd1358,-16'd1716,16'd144,16'd3164,16'd7773,-16'd7686};
dout[540]={ 16'd5317,-16'd1979,16'd5173,-16'd2875,-16'd3765,16'd4287,16'd1332,-16'd5020,16'd2903,16'd4074,16'd5785,16'd31,16'd2550,-16'd10895,16'd4842,16'd6582,-16'd607,-16'd1198,16'd2783,16'd649,-16'd4044,-16'd4528,-16'd10019,-16'd3213,16'd11523,-16'd4516,16'd1813,16'd2966,-16'd3204,16'd5502,-16'd7195,-16'd1293,16'd4405,-16'd7058,16'd11070,16'd2700};
dout[541]={ 16'd4993,16'd2780,-16'd714,-16'd7592,16'd6180,16'd5828,16'd2217,-16'd371,-16'd1967,16'd7954,16'd4533,-16'd5966,-16'd4600,-16'd3654,-16'd1048,16'd929,-16'd7173,16'd2993,16'd615,-16'd7092,-16'd6649,-16'd1089,-16'd329,-16'd4742,-16'd3379,16'd1598,-16'd1368,16'd5568,-16'd4046,16'd31,16'd295,-16'd959,16'd1142,-16'd6783,-16'd5790,16'd6175};
dout[542]={ -16'd4475,16'd4670,-16'd3855,-16'd3891,-16'd9117,-16'd2629,16'd2401,-16'd6560,-16'd2516,16'd6483,-16'd5837,-16'd11849,16'd1861,-16'd93,-16'd4324,16'd659,-16'd1241,16'd5465,-16'd1705,16'd6367,-16'd8165,-16'd2868,-16'd156,-16'd7969,-16'd2971,-16'd1054,-16'd9582,16'd6099,16'd2002,-16'd1687,-16'd6821,16'd2460,16'd741,-16'd902,-16'd5965,16'd4297};
dout[543]={ 16'd4838,-16'd705,16'd1424,-16'd4413,-16'd5146,-16'd5564,-16'd6968,-16'd978,-16'd4175,16'd9388,-16'd5437,16'd3573,16'd6827,-16'd451,16'd218,16'd3003,16'd4516,-16'd9554,-16'd386,-16'd629,16'd4833,-16'd9547,16'd208,-16'd9062,16'd6038,16'd5801,16'd2993,16'd3522,-16'd4100,-16'd2004,16'd5530,16'd5302,16'd8706,16'd2154,16'd3082,-16'd5857};
dout[544]={ 16'd5167,16'd3928,16'd699,16'd6034,-16'd6758,-16'd6458,16'd5798,-16'd6425,16'd3826,-16'd5688,-16'd10934,-16'd340,-16'd8053,-16'd3646,16'd4437,16'd4924,16'd1615,-16'd11491,16'd4019,-16'd1157,16'd6646,-16'd2282,-16'd2061,16'd3852,-16'd1004,-16'd5268,-16'd3111,16'd7144,16'd7771,16'd746,16'd5487,16'd4162,16'd5292,16'd9095,16'd1750,16'd5638};
dout[545]={ 16'd7127,-16'd768,-16'd5386,-16'd3764,-16'd4003,-16'd819,16'd4082,16'd3147,-16'd7133,-16'd5322,-16'd2257,-16'd2729,-16'd387,16'd5309,16'd3194,-16'd2096,16'd2400,-16'd3070,16'd1345,16'd6310,16'd3445,16'd2399,16'd4617,16'd1479,16'd3001,-16'd4658,-16'd7018,-16'd7939,16'd2627,16'd5510,-16'd583,-16'd2320,16'd3559,16'd3111,16'd1884,-16'd3474};
dout[546]={ 16'd4038,16'd4342,16'd4362,16'd5620,-16'd8755,16'd4414,16'd6357,-16'd2955,-16'd895,-16'd4146,-16'd4251,-16'd3198,-16'd8352,-16'd7056,-16'd1420,16'd2906,16'd1638,-16'd1303,-16'd5273,16'd4501,16'd6860,-16'd1826,-16'd654,16'd5717,-16'd2361,16'd747,16'd1826,16'd2058,-16'd7146,-16'd1910,-16'd7280,16'd6202,16'd3758,16'd7050,-16'd1688,-16'd574};
dout[547]={ -16'd707,-16'd6909,16'd2701,-16'd3553,-16'd1281,16'd5724,16'd2464,16'd3504,16'd5241,16'd2332,16'd3555,-16'd1596,-16'd6673,16'd2414,-16'd4040,-16'd6388,-16'd4652,16'd8,-16'd2019,16'd2715,16'd4975,-16'd710,16'd4101,16'd1825,16'd1389,-16'd6575,16'd6439,16'd1998,16'd2169,16'd4329,16'd3521,-16'd3173,16'd3660,-16'd3640,-16'd2801,16'd7659};
dout[548]={ -16'd6857,-16'd1875,16'd5694,16'd4961,-16'd7983,-16'd3363,16'd2001,16'd1239,16'd2249,16'd4550,-16'd1480,-16'd7357,-16'd4552,16'd3820,16'd250,-16'd2978,16'd115,-16'd1822,-16'd1802,-16'd1071,16'd157,16'd7255,16'd426,-16'd1540,16'd2957,-16'd6834,16'd3160,-16'd672,16'd6047,16'd2053,-16'd5832,-16'd3791,-16'd7490,-16'd3807,-16'd448,16'd8185};
dout[549]={ 16'd23,-16'd2297,-16'd4367,-16'd1739,-16'd4241,16'd2178,-16'd7921,16'd4116,-16'd3320,-16'd2175,-16'd654,-16'd2660,-16'd6424,16'd2516,16'd4608,16'd3801,-16'd5890,16'd2507,-16'd6780,16'd4111,-16'd634,-16'd6047,16'd5408,16'd2529,16'd4533,16'd2141,-16'd5907,16'd2114,-16'd3699,-16'd2467,16'd3236,-16'd3158,-16'd1617,-16'd1929,-16'd3171,-16'd6481};
dout[550]={ -16'd2354,-16'd1742,16'd3001,16'd9574,-16'd7863,-16'd7634,16'd653,16'd1711,16'd2401,16'd6127,16'd6529,-16'd3528,-16'd1224,-16'd3508,-16'd8234,16'd11511,-16'd2799,16'd261,-16'd4913,-16'd6588,16'd5808,-16'd6860,-16'd8295,16'd5956,16'd827,-16'd488,16'd5198,-16'd1005,-16'd4362,-16'd1858,-16'd6655,16'd8603,16'd2120,16'd5331,16'd4184,16'd4336};
dout[551]={ 16'd5076,-16'd4974,-16'd5058,-16'd5870,16'd4254,-16'd1150,-16'd8019,-16'd2061,-16'd71,16'd1263,16'd2786,-16'd6224,-16'd3375,16'd3569,-16'd9042,-16'd5617,16'd4618,16'd913,-16'd7552,-16'd4432,16'd6771,-16'd8041,-16'd6738,16'd250,-16'd500,-16'd2016,-16'd9561,-16'd5355,16'd1353,16'd497,16'd4697,-16'd4596,16'd4443,-16'd341,-16'd1342,16'd1547};
dout[552]={ 16'd1502,-16'd897,-16'd10828,-16'd10211,-16'd3580,16'd8957,-16'd4504,16'd4142,-16'd2795,16'd10261,16'd1152,-16'd10959,16'd5208,-16'd26,-16'd9841,-16'd9351,16'd4227,16'd2943,16'd2085,-16'd6201,-16'd2101,-16'd1096,-16'd938,16'd2380,16'd8135,-16'd1815,16'd2243,16'd3388,-16'd10076,16'd3642,-16'd1195,16'd3101,16'd1115,-16'd489,-16'd881,16'd224};
dout[553]={ 16'd2405,16'd6412,-16'd6407,-16'd295,-16'd4306,-16'd6200,-16'd4004,16'd1855,-16'd7089,-16'd4704,-16'd11535,-16'd9932,16'd2717,-16'd1333,-16'd4749,-16'd2238,16'd4497,-16'd11144,16'd866,16'd2866,16'd5118,-16'd2384,-16'd101,-16'd7299,-16'd6296,16'd3239,16'd4162,16'd2716,-16'd5685,16'd3919,16'd1294,16'd2000,-16'd2814,16'd7373,-16'd5985,-16'd1674};
dout[554]={ 16'd4516,16'd2311,16'd3378,16'd3762,16'd6069,-16'd807,16'd1087,16'd5554,16'd3980,-16'd3940,-16'd6939,-16'd4702,-16'd1768,16'd7085,16'd7794,16'd2812,-16'd2737,-16'd4435,-16'd8096,-16'd817,-16'd1033,16'd6357,16'd2112,-16'd2773,16'd618,16'd2402,16'd7823,16'd401,16'd280,-16'd1492,-16'd7732,-16'd4653,-16'd3518,16'd7411,-16'd3035,16'd4040};
dout[555]={ -16'd2347,-16'd1388,16'd3194,16'd5767,-16'd4960,16'd7556,16'd1032,-16'd3143,16'd6432,-16'd770,16'd4428,16'd3842,16'd3181,16'd7430,16'd2631,-16'd4766,-16'd7580,-16'd4756,-16'd6900,16'd2376,16'd1645,16'd2552,16'd5662,16'd4872,-16'd4972,16'd2321,16'd3281,16'd303,16'd7435,16'd4158,-16'd1762,16'd8400,16'd5782,16'd6396,-16'd3825,16'd6396};
dout[556]={ -16'd6279,16'd2768,-16'd5687,-16'd2902,-16'd3472,-16'd1056,-16'd5585,16'd4323,-16'd3027,16'd2048,-16'd2059,-16'd2178,-16'd5045,16'd3129,-16'd4412,-16'd3972,16'd2267,-16'd5917,16'd3850,-16'd6091,-16'd5472,-16'd6792,-16'd3370,16'd1071,16'd5537,-16'd4880,-16'd3432,-16'd2052,16'd3417,16'd4382,16'd1927,16'd4634,16'd6112,16'd4207,16'd3129,16'd1517};
dout[557]={ 16'd1713,16'd5217,-16'd1077,-16'd3687,-16'd5038,-16'd3612,-16'd4737,16'd935,16'd2196,16'd5091,16'd6235,16'd1873,-16'd56,-16'd221,-16'd2681,-16'd1238,-16'd5035,-16'd3541,16'd6483,-16'd3282,-16'd6389,16'd2528,16'd1629,-16'd531,16'd5760,-16'd2671,-16'd3525,-16'd5436,16'd4679,16'd2094,-16'd2330,-16'd816,-16'd5934,16'd4282,-16'd1789,16'd1257};
dout[558]={ 16'd3845,16'd3346,16'd599,16'd2926,-16'd2040,-16'd3294,16'd1343,16'd5100,16'd4122,-16'd6243,-16'd2135,16'd6298,-16'd6271,-16'd1198,-16'd5868,-16'd5072,16'd4757,-16'd7137,-16'd4559,-16'd120,-16'd110,-16'd603,-16'd1254,16'd3863,16'd4941,-16'd6515,16'd5695,-16'd4823,16'd4578,-16'd427,-16'd6329,16'd3943,-16'd2715,-16'd7603,16'd3837,-16'd4018};
dout[559]={ 16'd1198,-16'd691,16'd357,-16'd5614,-16'd4100,-16'd976,-16'd5717,-16'd6251,-16'd6877,-16'd5293,16'd3281,16'd2633,16'd6812,-16'd3,-16'd133,16'd4778,-16'd1437,-16'd2328,16'd4984,-16'd7471,-16'd4731,-16'd591,-16'd4691,16'd1477,-16'd7286,16'd2933,16'd4573,16'd2228,-16'd1260,16'd4062,16'd6955,16'd3975,16'd4789,-16'd5370,-16'd6612,16'd1771};
dout[560]={ 16'd757,-16'd319,-16'd1350,16'd5498,-16'd4583,-16'd8335,16'd5262,-16'd4881,16'd3370,16'd2053,16'd546,16'd6347,16'd8443,-16'd10976,16'd4580,-16'd2658,-16'd5762,-16'd2591,16'd262,-16'd8171,16'd177,-16'd4005,-16'd7183,-16'd5046,16'd576,-16'd2623,16'd5829,16'd6965,16'd2615,16'd1468,-16'd8168,-16'd977,16'd5177,-16'd5375,16'd746,16'd2901};
dout[561]={ -16'd316,-16'd3731,-16'd4530,16'd32,-16'd3026,-16'd523,16'd3303,-16'd5880,16'd1637,16'd5932,-16'd5035,16'd3528,16'd488,-16'd10359,-16'd7965,16'd731,16'd366,16'd1108,-16'd53,16'd6064,16'd4881,-16'd2827,16'd1192,-16'd67,-16'd1605,-16'd3250,-16'd9965,16'd2524,-16'd8290,-16'd3564,16'd4726,-16'd321,16'd5225,-16'd9017,16'd6468,16'd5527};
dout[562]={ 16'd1635,-16'd7271,-16'd9017,-16'd4705,16'd3322,-16'd1010,16'd2083,-16'd664,-16'd1926,16'd4303,-16'd5069,16'd1693,-16'd6029,16'd3608,16'd66,-16'd8135,16'd4757,-16'd5324,-16'd72,16'd1538,-16'd4683,-16'd1756,-16'd5805,-16'd5378,16'd7271,-16'd3205,16'd2545,-16'd2604,-16'd8939,16'd5285,-16'd7636,16'd5302,-16'd4166,-16'd11963,-16'd4415,16'd3117};
dout[563]={ -16'd2592,16'd3686,-16'd6783,-16'd6762,16'd6243,16'd8186,-16'd6630,-16'd4742,-16'd3123,-16'd8150,16'd828,-16'd6299,16'd2606,-16'd251,-16'd1620,-16'd3522,16'd2217,16'd2390,-16'd439,16'd677,-16'd5941,16'd2175,16'd3851,-16'd6669,16'd1685,-16'd4124,-16'd5765,-16'd1539,-16'd4992,-16'd1534,-16'd3333,16'd1794,16'd7754,16'd322,-16'd1275,16'd848};
dout[564]={ 16'd4278,16'd3425,16'd6190,16'd7750,-16'd2391,16'd4613,-16'd8296,-16'd3551,16'd1330,-16'd7662,-16'd4953,-16'd3928,-16'd2977,-16'd1882,-16'd2171,-16'd6856,-16'd1517,16'd1824,16'd2717,-16'd5772,16'd6398,16'd6877,-16'd705,-16'd7228,-16'd142,-16'd388,-16'd1810,16'd4452,-16'd107,-16'd8031,-16'd6270,16'd2884,-16'd882,16'd7550,-16'd4603,16'd5621};
dout[565]={ 16'd34,-16'd1711,16'd5720,-16'd1974,-16'd6584,16'd3569,-16'd2936,-16'd4174,-16'd3490,16'd697,16'd1648,-16'd1237,16'd5487,-16'd755,16'd2578,16'd3934,-16'd3,-16'd2678,16'd2895,-16'd4214,16'd2630,-16'd7078,-16'd1549,-16'd5460,16'd2275,16'd6326,16'd16,-16'd6673,16'd7469,16'd484,16'd827,-16'd2370,16'd917,16'd4399,-16'd8057,16'd5252};
dout[566]={ 16'd6713,-16'd1777,-16'd164,16'd4557,-16'd5003,-16'd4047,16'd3100,-16'd4181,-16'd3111,-16'd4827,16'd1477,16'd1962,-16'd5196,-16'd3439,16'd6976,-16'd7294,16'd5515,-16'd5811,16'd4928,-16'd4600,16'd7131,-16'd7201,-16'd530,16'd816,-16'd6691,16'd4314,16'd2789,16'd7613,16'd6446,16'd3439,-16'd5493,-16'd3081,-16'd2957,-16'd4731,-16'd1659,16'd4293};
dout[567]={ -16'd3467,-16'd5871,16'd39,16'd7804,-16'd7358,-16'd2452,-16'd5919,-16'd7786,16'd1072,16'd287,-16'd3877,16'd6827,-16'd5975,-16'd4099,16'd1270,16'd580,-16'd1200,-16'd4154,16'd5249,16'd936,16'd5730,-16'd7534,-16'd394,-16'd2865,16'd3233,16'd1153,-16'd499,16'd1183,16'd3931,16'd919,16'd1754,-16'd5370,-16'd750,-16'd3117,16'd4725,16'd1400};
dout[568]={ -16'd7089,16'd5045,16'd7024,16'd3709,16'd1789,-16'd2563,16'd6228,16'd5241,-16'd7716,-16'd5878,-16'd767,-16'd7175,-16'd3476,16'd4072,-16'd2780,-16'd3743,16'd5041,-16'd3471,-16'd3867,-16'd825,-16'd246,16'd4064,-16'd397,-16'd7444,16'd3398,16'd1729,-16'd845,16'd3484,-16'd4699,16'd1449,-16'd5392,16'd5714,-16'd345,-16'd6709,-16'd4547,16'd4819};
dout[569]={ 16'd1768,-16'd6686,16'd5775,16'd7258,16'd1053,-16'd2566,16'd72,16'd6092,-16'd8685,-16'd643,-16'd3478,16'd2476,16'd4200,16'd4632,16'd2549,16'd2400,-16'd3998,16'd1569,16'd4549,-16'd2133,-16'd2989,-16'd8252,16'd6135,16'd6998,16'd2463,-16'd882,-16'd782,16'd5446,-16'd7043,-16'd1357,16'd2847,-16'd1892,16'd6901,16'd2627,16'd3941,-16'd353};
dout[570]={ -16'd4373,-16'd7147,16'd192,-16'd821,-16'd5624,-16'd8101,16'd1396,16'd6409,16'd4858,-16'd2471,-16'd833,-16'd6144,-16'd1510,-16'd5914,16'd1990,16'd2522,16'd4191,-16'd1084,16'd986,16'd1607,-16'd7296,-16'd5663,-16'd487,-16'd4191,-16'd1827,16'd1407,-16'd3015,-16'd3634,-16'd7258,16'd4913,-16'd6868,16'd2011,16'd1250,-16'd6062,16'd6375,16'd1148};
dout[571]={ 16'd1871,16'd4092,-16'd9147,-16'd2526,16'd4530,-16'd2785,16'd1298,-16'd5129,-16'd752,-16'd6791,-16'd3245,-16'd9444,16'd4387,-16'd3978,-16'd3809,-16'd4959,-16'd9245,-16'd1800,16'd4376,16'd6522,16'd4009,16'd2245,16'd5351,16'd34,16'd9009,16'd7982,-16'd7410,16'd2406,16'd4564,-16'd2203,-16'd2826,16'd3708,16'd4232,-16'd8132,-16'd1997,-16'd3307};
dout[572]={ -16'd3454,16'd2220,-16'd2434,16'd4168,-16'd129,16'd5512,16'd5542,-16'd8152,-16'd2161,16'd1685,-16'd603,-16'd1077,16'd5618,-16'd3870,-16'd2320,-16'd10591,-16'd4960,-16'd2275,-16'd8934,16'd1167,-16'd2353,-16'd1213,-16'd3157,-16'd8400,-16'd2360,-16'd5618,-16'd6607,-16'd4462,16'd2143,16'd79,16'd4010,16'd4439,16'd7175,-16'd10836,16'd10934,-16'd874};
dout[573]={ 16'd130,16'd3960,-16'd8242,-16'd6177,-16'd2966,16'd231,16'd3702,-16'd1487,-16'd6203,-16'd9716,-16'd5913,-16'd1033,16'd5259,16'd4088,-16'd2997,-16'd8568,-16'd7012,-16'd7138,16'd4620,16'd3923,-16'd1732,-16'd4371,16'd204,-16'd1579,-16'd4533,16'd364,-16'd4188,16'd1363,16'd7069,-16'd5364,16'd2795,-16'd1691,-16'd4432,16'd116,16'd3843,16'd2760};
dout[574]={ -16'd1025,-16'd839,-16'd7875,16'd1710,-16'd3194,16'd2157,16'd3101,16'd1219,-16'd5807,-16'd6719,16'd3463,16'd1606,-16'd795,16'd1764,16'd2361,-16'd4266,-16'd3843,16'd1012,16'd5535,-16'd596,16'd1272,16'd1200,16'd7443,-16'd3168,16'd534,-16'd229,16'd6538,-16'd5879,-16'd618,-16'd5429,-16'd7983,16'd2170,-16'd7207,-16'd6123,16'd2017,16'd7418};
dout[575]={ -16'd2093,-16'd6764,-16'd2156,-16'd4012,-16'd7361,16'd736,-16'd3592,-16'd1059,-16'd471,-16'd2583,16'd2341,16'd217,16'd4290,-16'd6305,-16'd2939,16'd2948,-16'd3072,-16'd3242,16'd5787,-16'd4251,16'd2771,16'd4247,-16'd3389,16'd3637,-16'd3683,-16'd7716,16'd1910,16'd6487,16'd4028,16'd5613,-16'd6117,-16'd3516,16'd5231,16'd9024,-16'd9830,-16'd6966};
dout[576]={ -16'd5416,16'd3978,16'd2759,-16'd1124,-16'd1671,-16'd2209,-16'd228,-16'd6179,16'd5624,-16'd968,-16'd1587,-16'd1863,-16'd2878,16'd3062,16'd6577,-16'd1828,-16'd1212,-16'd284,-16'd6523,16'd3975,-16'd7619,-16'd4126,-16'd1047,-16'd2183,-16'd5663,16'd5297,-16'd7609,16'd2197,-16'd3140,-16'd3061,-16'd4957,16'd120,-16'd4717,16'd2027,-16'd1515,-16'd3477};
dout[577]={ -16'd4441,-16'd529,16'd4703,16'd5374,16'd6330,-16'd5093,16'd2959,16'd4325,-16'd3128,-16'd5884,16'd1541,-16'd3812,-16'd5958,-16'd3410,16'd248,-16'd3254,16'd339,16'd3242,16'd3544,16'd2249,16'd3302,16'd2360,16'd314,-16'd6148,-16'd4882,-16'd8493,-16'd204,16'd1605,-16'd8700,16'd5570,-16'd6817,-16'd4814,16'd2423,16'd17,-16'd3126,-16'd5110};
dout[578]={ -16'd5029,-16'd3499,16'd3327,-16'd5403,16'd4696,16'd3444,-16'd5302,-16'd3379,16'd5059,-16'd3361,-16'd3951,16'd5725,-16'd9,16'd2230,-16'd4368,-16'd332,-16'd4299,16'd3915,16'd2218,-16'd4351,16'd5314,-16'd6529,16'd2939,-16'd1637,16'd1139,-16'd2560,-16'd418,16'd5099,16'd2957,16'd4759,16'd4335,-16'd5149,16'd8684,16'd4426,-16'd1470,16'd6827};
dout[579]={ -16'd7265,16'd5394,-16'd6,16'd4815,16'd396,16'd6836,-16'd6412,16'd3153,16'd4719,16'd94,16'd5281,-16'd5087,-16'd925,16'd2735,16'd2061,16'd3600,16'd3263,-16'd8849,-16'd393,-16'd1214,16'd5935,16'd4381,-16'd3558,16'd3538,-16'd145,-16'd3951,16'd5183,-16'd1133,-16'd1681,-16'd2379,-16'd2625,-16'd4821,-16'd4517,16'd2256,-16'd256,16'd5147};
dout[580]={ 16'd3835,-16'd11579,-16'd7410,16'd4267,16'd4846,-16'd1499,16'd1456,-16'd1482,-16'd6819,16'd3357,16'd3427,-16'd3616,-16'd6153,16'd1330,-16'd6130,-16'd3203,-16'd254,16'd4427,16'd6488,-16'd3297,-16'd5947,-16'd239,16'd6304,-16'd1498,16'd4413,16'd2417,16'd3961,16'd6437,16'd5275,-16'd1335,-16'd4351,16'd3946,-16'd1021,-16'd5785,16'd5606,16'd2506};
dout[581]={ -16'd401,-16'd3631,-16'd5469,-16'd2914,-16'd4454,-16'd5522,-16'd6659,16'd3172,16'd1003,-16'd4984,-16'd6477,-16'd2266,16'd3796,16'd4895,-16'd3864,16'd4523,-16'd131,16'd1839,16'd6363,16'd1324,-16'd4788,-16'd3693,-16'd1774,16'd6709,-16'd4470,-16'd3144,16'd4600,-16'd5308,-16'd7886,16'd6816,16'd2710,-16'd317,-16'd3034,-16'd4839,16'd1566,-16'd8931};
dout[582]={ 16'd3359,-16'd2372,-16'd4408,-16'd9990,-16'd2750,16'd6939,-16'd337,16'd4754,-16'd3752,16'd7089,16'd4357,16'd2319,-16'd642,16'd1258,-16'd5871,-16'd8026,-16'd7740,-16'd4559,16'd2272,16'd5885,-16'd363,-16'd4640,16'd1213,-16'd3884,16'd5547,16'd2414,-16'd132,16'd3513,16'd5220,16'd9375,16'd1356,16'd6849,16'd3665,-16'd776,16'd6484,-16'd2826};
dout[583]={ -16'd3135,16'd4068,-16'd7717,-16'd2509,-16'd5350,16'd4722,-16'd5552,-16'd2134,16'd4641,-16'd3994,-16'd5243,-16'd3033,16'd7113,-16'd330,16'd3901,-16'd1754,16'd6140,-16'd3540,-16'd6496,16'd2976,16'd5973,-16'd4081,-16'd4251,16'd6307,16'd2531,16'd4424,16'd1023,16'd5281,16'd7567,16'd2618,-16'd3698,-16'd6959,16'd1015,16'd652,16'd1137,16'd7335};
dout[584]={ 16'd1298,16'd1463,-16'd459,-16'd3883,16'd2564,-16'd3506,16'd3239,16'd2810,-16'd1618,-16'd7069,-16'd4808,16'd4683,16'd6614,16'd6257,16'd1671,16'd983,16'd3347,16'd2591,-16'd719,-16'd6731,16'd5296,16'd4282,16'd711,-16'd4042,-16'd6747,-16'd3913,-16'd2424,16'd2523,16'd2275,-16'd2794,16'd4822,-16'd9585,-16'd5568,16'd3211,-16'd3027,16'd5065};
dout[585]={ -16'd6362,16'd3047,16'd7143,-16'd1773,-16'd3754,16'd6387,16'd20,-16'd4503,-16'd8069,16'd1292,16'd3060,-16'd3596,16'd4979,16'd136,16'd2620,-16'd4302,16'd4041,16'd4194,16'd7231,-16'd178,16'd5050,16'd5058,-16'd2345,-16'd5205,16'd6741,16'd1833,16'd4579,-16'd2119,-16'd5520,16'd345,16'd5210,16'd4832,16'd6590,-16'd3242,16'd1728,16'd1561};
dout[586]={ -16'd1313,16'd3561,-16'd2352,16'd7611,-16'd1380,-16'd6129,-16'd6055,16'd4533,16'd3651,-16'd1409,16'd754,-16'd33,16'd5800,16'd8218,-16'd329,16'd4288,16'd3748,-16'd1648,16'd3213,-16'd1633,-16'd7692,-16'd5878,16'd57,-16'd5214,-16'd3518,-16'd6884,16'd5885,-16'd3295,-16'd247,16'd371,16'd671,-16'd4331,16'd548,16'd1965,-16'd3612,16'd7264};
dout[587]={ -16'd2481,16'd539,-16'd3997,16'd8729,-16'd4425,-16'd1292,-16'd3349,-16'd5183,16'd2996,-16'd4091,-16'd2309,16'd1076,-16'd452,16'd3596,-16'd1308,-16'd2669,-16'd8089,-16'd4653,16'd3271,16'd5645,-16'd4291,16'd1971,16'd4706,16'd5284,-16'd4101,-16'd1289,-16'd5535,-16'd514,16'd1474,16'd1776,16'd4968,16'd894,16'd2262,-16'd3447,-16'd5837,16'd3805};
dout[588]={ -16'd6447,16'd3695,16'd1523,16'd4760,16'd1408,-16'd5609,-16'd4818,-16'd5019,16'd3939,-16'd3834,16'd4630,-16'd1538,-16'd6329,-16'd5624,16'd3567,16'd2167,16'd3933,16'd2857,-16'd2432,16'd5039,16'd1259,16'd5309,-16'd4130,16'd4473,16'd3210,16'd3118,16'd6032,-16'd3528,16'd923,16'd1412,-16'd4487,-16'd2651,-16'd1203,-16'd4654,-16'd4027,16'd7089};
dout[589]={ -16'd889,-16'd5427,16'd589,16'd3550,16'd3724,16'd2757,16'd5612,-16'd2030,-16'd4129,16'd92,-16'd723,16'd6859,-16'd3124,16'd30,-16'd3106,16'd1687,16'd3166,16'd4817,-16'd4511,-16'd567,16'd3468,16'd29,-16'd534,16'd5958,-16'd5143,-16'd33,-16'd7454,16'd6179,16'd748,16'd6516,16'd5935,16'd4283,-16'd4354,16'd4331,16'd703,-16'd6045};
dout[590]={ -16'd12003,16'd3056,16'd988,16'd2057,-16'd371,-16'd2450,16'd546,-16'd987,16'd4850,-16'd3067,-16'd1698,-16'd1195,-16'd2844,16'd2679,16'd3836,-16'd9408,-16'd9799,-16'd2413,-16'd4123,-16'd5757,16'd5068,16'd3770,16'd3124,-16'd6389,16'd4434,16'd7584,-16'd5149,16'd628,16'd3251,-16'd3169,16'd5236,16'd5637,16'd11927,-16'd2125,16'd338,-16'd7426};
dout[591]={ -16'd2150,16'd3269,-16'd1043,16'd895,16'd2085,-16'd2099,16'd4618,-16'd1591,-16'd8863,16'd5326,-16'd3999,-16'd9386,-16'd1949,16'd3350,16'd1947,-16'd493,-16'd1770,-16'd10,-16'd5344,16'd8022,-16'd8370,-16'd483,16'd4897,-16'd1022,-16'd7422,16'd2813,-16'd6521,16'd7784,-16'd5727,16'd6190,16'd1884,16'd2597,16'd4411,-16'd7311,16'd2882,-16'd538};
dout[592]={ -16'd8719,16'd5517,-16'd7607,-16'd8063,16'd7103,16'd5368,-16'd4924,16'd4424,-16'd7686,16'd142,16'd5514,-16'd2032,-16'd7245,16'd3852,-16'd6487,-16'd3997,16'd4737,-16'd6750,16'd3359,-16'd5925,16'd5542,-16'd6925,16'd2985,-16'd8897,-16'd2558,16'd6229,-16'd6522,16'd1093,16'd8308,16'd7724,16'd1848,-16'd5613,16'd1840,-16'd8413,-16'd1877,16'd396};
dout[593]={ -16'd3027,-16'd5480,16'd2803,-16'd2199,-16'd3540,16'd21,-16'd2352,-16'd3984,-16'd5088,-16'd504,-16'd544,16'd3292,16'd2296,-16'd6838,16'd6300,-16'd12742,-16'd4034,-16'd4252,-16'd4410,-16'd4499,-16'd1802,-16'd3868,16'd6015,-16'd3477,-16'd4592,-16'd209,-16'd2998,-16'd212,16'd1402,-16'd1798,-16'd603,-16'd5510,-16'd5350,16'd5108,-16'd4632,-16'd6300};
dout[594]={ 16'd3810,-16'd559,-16'd955,16'd3698,-16'd6972,-16'd3263,16'd2799,-16'd3163,-16'd2658,-16'd4339,16'd5422,-16'd7254,-16'd7352,-16'd326,-16'd1699,-16'd3651,-16'd5196,-16'd6845,16'd3406,16'd1258,-16'd4590,-16'd2628,-16'd4400,16'd364,16'd2701,-16'd4113,16'd8190,-16'd8269,16'd238,-16'd1267,-16'd1927,16'd4831,-16'd6720,-16'd3752,-16'd11440,16'd118};
dout[595]={ 16'd820,16'd5142,16'd5183,16'd8126,-16'd6767,-16'd1228,16'd7019,-16'd3191,-16'd3277,-16'd5204,16'd4103,-16'd8071,16'd5938,-16'd1009,-16'd1538,16'd2452,16'd4263,-16'd2554,-16'd2862,16'd2635,-16'd1963,-16'd117,-16'd4299,16'd1501,16'd2470,-16'd2759,-16'd2959,16'd5186,-16'd6372,-16'd2341,16'd1697,-16'd4074,16'd4997,16'd8189,-16'd5517,-16'd2038};
dout[596]={ 16'd314,-16'd4419,16'd890,-16'd1988,-16'd3785,-16'd6493,-16'd4246,16'd2551,16'd4808,16'd2925,16'd3290,-16'd5725,16'd6268,16'd6361,-16'd1196,-16'd8249,16'd4437,-16'd268,16'd7056,-16'd1192,16'd4474,-16'd4452,16'd883,-16'd2038,-16'd3670,-16'd263,-16'd4724,-16'd7320,16'd3026,16'd1546,-16'd2374,16'd4003,16'd9038,-16'd3063,-16'd4839,16'd3482};
dout[597]={ -16'd3554,-16'd3733,-16'd383,-16'd2217,16'd4246,-16'd3151,16'd2739,-16'd1004,16'd1620,-16'd4148,16'd3956,-16'd794,16'd3333,-16'd143,16'd7011,16'd5989,-16'd286,16'd4700,-16'd2769,-16'd4030,-16'd7809,-16'd3180,-16'd8697,-16'd6754,-16'd8254,-16'd5508,16'd147,-16'd1980,-16'd5947,16'd4258,16'd3558,16'd5079,-16'd4448,16'd8159,-16'd8134,-16'd6453};
dout[598]={ 16'd2343,-16'd5622,-16'd2804,-16'd601,16'd4879,-16'd1421,16'd3389,-16'd641,-16'd3576,16'd1999,-16'd6281,16'd5040,16'd2621,16'd2924,16'd3098,16'd3506,16'd4204,16'd661,-16'd6631,16'd3110,16'd2515,16'd2552,16'd6511,16'd5802,-16'd6501,-16'd5065,-16'd1726,16'd5158,-16'd318,-16'd5646,-16'd2281,-16'd3019,16'd4006,16'd5282,16'd4165,16'd1181};
dout[599]={ 16'd1170,-16'd2309,16'd7416,16'd4839,-16'd4636,16'd7177,-16'd1570,16'd7578,16'd4333,16'd6609,-16'd4532,-16'd2047,-16'd2078,16'd1098,-16'd4492,16'd1007,16'd401,-16'd5724,16'd3943,16'd5552,-16'd1116,-16'd3035,16'd221,-16'd8051,-16'd1464,-16'd5853,-16'd802,16'd4313,-16'd6354,-16'd3620,-16'd2928,-16'd2870,-16'd4363,16'd1844,16'd3286,-16'd3931};
dout[600]={ -16'd4854,-16'd818,-16'd475,-16'd2540,16'd37,16'd3265,16'd6465,-16'd2995,16'd4163,16'd7374,-16'd10789,-16'd3914,-16'd1802,16'd3000,-16'd5116,16'd2667,-16'd3379,-16'd464,-16'd7409,-16'd1841,-16'd7979,-16'd9474,-16'd1045,-16'd765,16'd2224,16'd1776,-16'd2383,16'd11993,16'd2545,-16'd1723,-16'd5066,-16'd9930,-16'd2274,-16'd7330,-16'd7479,16'd5231};
dout[601]={ -16'd902,16'd5386,16'd8035,16'd1468,16'd2073,-16'd6353,16'd6601,-16'd1910,-16'd2634,-16'd5190,-16'd3265,-16'd1662,16'd6060,-16'd2515,16'd4767,16'd5180,-16'd5209,-16'd8735,-16'd3315,-16'd814,-16'd9770,-16'd3231,-16'd7791,16'd1033,16'd3137,16'd137,16'd8366,-16'd2708,-16'd9823,16'd1317,16'd3960,-16'd1200,16'd3884,-16'd1864,16'd4434,16'd3476};
dout[602]={ -16'd3835,-16'd1460,16'd862,-16'd1042,-16'd4920,-16'd6084,-16'd1695,-16'd2052,-16'd5252,16'd8509,-16'd10820,-16'd1930,-16'd2117,-16'd7325,-16'd232,-16'd5877,16'd1740,16'd6138,-16'd3016,16'd2918,16'd3102,-16'd1864,16'd4725,16'd1337,-16'd7592,16'd5703,16'd4719,16'd2509,-16'd4309,-16'd4283,16'd5960,16'd1776,-16'd4750,16'd565,16'd6973,16'd5198};
dout[603]={ -16'd3945,16'd3483,-16'd569,16'd5538,-16'd1531,16'd4517,16'd2297,-16'd6373,-16'd5142,16'd5802,-16'd6605,16'd1534,-16'd5855,16'd3372,-16'd1752,-16'd5715,-16'd7275,-16'd4034,16'd4663,-16'd1783,16'd4180,-16'd5175,16'd4479,-16'd9249,16'd5665,-16'd1881,16'd4507,16'd7379,16'd687,16'd1643,16'd3201,16'd1339,-16'd3175,16'd5092,16'd3497,16'd5967};
dout[604]={ 16'd4690,16'd8121,16'd9516,16'd5500,-16'd3548,16'd6459,-16'd7004,-16'd7515,-16'd5397,16'd3256,-16'd2398,-16'd3876,16'd1599,-16'd5406,16'd2974,16'd5313,-16'd4854,16'd1616,16'd6542,-16'd2040,-16'd4737,16'd3390,-16'd4503,-16'd3961,-16'd3480,16'd1194,16'd7679,16'd4334,-16'd8244,16'd9095,-16'd5649,-16'd2578,-16'd585,16'd4698,-16'd7734,16'd1243};
dout[605]={ 16'd32,16'd403,16'd2394,16'd2634,16'd2594,-16'd6252,16'd3304,16'd4260,-16'd4751,-16'd3297,16'd2275,16'd101,-16'd3551,16'd1360,16'd4818,-16'd157,16'd4069,16'd2822,-16'd4941,-16'd3954,16'd4397,16'd3452,-16'd1126,16'd2534,-16'd7362,16'd5489,-16'd4946,16'd4391,16'd3464,-16'd3323,16'd4749,16'd5076,16'd5602,16'd1217,16'd2466,16'd2205};
dout[606]={ 16'd1804,-16'd442,-16'd1979,16'd3716,16'd7695,16'd689,16'd3051,16'd5985,-16'd292,16'd6945,16'd438,16'd7139,-16'd1482,-16'd2584,-16'd916,16'd162,16'd1029,16'd4935,16'd7748,16'd5510,-16'd4975,-16'd4590,16'd5437,-16'd1589,-16'd5173,-16'd2495,-16'd6193,-16'd4813,-16'd367,16'd5341,16'd342,16'd4151,-16'd2670,16'd1072,16'd5650,-16'd2156};
dout[607]={ 16'd3818,-16'd6268,-16'd969,-16'd225,-16'd3264,-16'd1877,-16'd2347,16'd6577,-16'd8273,-16'd6713,-16'd6562,-16'd368,16'd5766,-16'd5578,-16'd3575,16'd6722,-16'd1438,16'd764,-16'd4653,-16'd919,16'd6496,-16'd7556,16'd986,-16'd1079,-16'd338,16'd727,16'd6231,-16'd7676,-16'd1305,16'd2066,16'd3820,16'd4052,16'd6288,16'd4970,16'd8033,-16'd553};
dout[608]={ 16'd1368,-16'd1903,16'd7233,16'd4689,-16'd3336,-16'd6740,16'd8008,16'd705,-16'd4929,16'd2435,16'd278,16'd4033,16'd5707,16'd4909,-16'd2147,16'd4826,-16'd3576,16'd728,16'd2458,-16'd576,-16'd493,-16'd3765,16'd2257,16'd319,-16'd3466,-16'd3751,16'd3001,-16'd1784,-16'd7471,16'd5521,-16'd2432,-16'd6373,-16'd2390,-16'd3617,-16'd88,-16'd6636};
dout[609]={ 16'd3666,16'd3927,-16'd3052,16'd1705,16'd1869,-16'd3587,-16'd2062,16'd5189,16'd843,16'd4329,-16'd41,-16'd5453,16'd4020,-16'd2760,16'd9144,-16'd3384,-16'd4396,-16'd6080,16'd6461,16'd2354,16'd3120,-16'd4100,16'd0,-16'd2181,16'd1430,16'd2657,16'd4244,-16'd6058,16'd5489,-16'd5496,16'd6886,16'd7065,-16'd5737,-16'd4912,16'd475,-16'd5773};
dout[610]={ 16'd4072,16'd4506,-16'd3918,16'd2069,-16'd7361,16'd2636,-16'd252,-16'd6819,16'd1588,16'd8466,-16'd8221,-16'd2134,16'd2271,-16'd3077,16'd4192,-16'd7770,-16'd2106,16'd143,-16'd6067,16'd279,-16'd28,16'd2691,-16'd3020,-16'd5150,-16'd1967,-16'd9773,16'd1882,16'd10316,-16'd1088,16'd4952,-16'd8964,-16'd2077,-16'd5058,16'd1436,16'd5044,-16'd7246};
dout[611]={ 16'd7125,-16'd626,16'd3817,-16'd9229,16'd4934,-16'd2240,-16'd2705,16'd1015,16'd1826,16'd2763,-16'd9249,16'd549,-16'd7687,-16'd5870,-16'd7918,-16'd2669,-16'd4142,16'd3794,16'd591,-16'd8671,-16'd522,16'd6232,-16'd1763,-16'd2710,16'd4963,-16'd8552,16'd4443,-16'd2601,-16'd501,16'd396,-16'd8238,16'd1696,16'd6237,-16'd5864,16'd103,16'd2177};
dout[612]={ 16'd5854,16'd1866,16'd207,16'd2226,16'd1629,-16'd4892,-16'd6426,-16'd741,16'd980,16'd342,-16'd8480,-16'd5186,-16'd1550,-16'd3698,-16'd5995,-16'd3545,16'd4927,16'd426,16'd4063,-16'd9592,-16'd70,-16'd3178,-16'd4658,16'd4010,-16'd7373,-16'd7502,-16'd464,-16'd4060,-16'd7317,-16'd4418,16'd2249,-16'd6721,-16'd7184,-16'd7821,16'd2535,-16'd6465};
dout[613]={ -16'd807,16'd9936,-16'd1539,-16'd1301,-16'd1586,16'd5934,16'd7272,16'd4266,16'd1421,-16'd2802,-16'd9161,-16'd1733,16'd5797,-16'd3188,16'd4218,-16'd5421,-16'd5947,16'd6640,16'd1518,16'd2803,-16'd7550,-16'd10287,-16'd2393,-16'd9844,16'd4012,16'd6224,-16'd5866,-16'd2867,16'd1072,-16'd3467,-16'd1276,-16'd3090,-16'd3548,16'd3129,-16'd6145,16'd776};
dout[614]={ 16'd5493,-16'd1823,16'd5621,-16'd2142,16'd5035,16'd3132,16'd2073,16'd3481,16'd1128,16'd1039,-16'd10656,16'd2852,16'd7129,-16'd6636,-16'd4096,16'd6213,16'd5166,-16'd3977,-16'd1598,-16'd3993,16'd6857,-16'd9637,-16'd1773,-16'd1505,-16'd470,16'd5673,16'd3343,16'd65,-16'd8016,-16'd4648,16'd2198,16'd8811,-16'd7707,16'd31,-16'd2722,16'd2392};
dout[615]={ 16'd39,-16'd2748,16'd4010,-16'd8338,-16'd4940,16'd3837,-16'd5928,-16'd8377,16'd5140,16'd1754,-16'd7929,16'd543,16'd2351,-16'd5608,-16'd5337,-16'd8606,16'd5381,16'd3391,-16'd2948,16'd3281,-16'd3091,-16'd1065,-16'd6525,-16'd7706,-16'd6741,-16'd3473,16'd277,16'd2981,16'd286,16'd5555,-16'd7742,-16'd3884,16'd2247,16'd3467,-16'd4619,16'd3495};
dout[616]={ 16'd2381,16'd1972,16'd5443,16'd4353,16'd6174,-16'd2096,-16'd4000,-16'd1474,16'd801,-16'd1784,16'd4011,16'd394,-16'd430,16'd1285,16'd2651,-16'd4709,16'd6664,16'd5770,16'd5393,16'd2767,16'd2721,-16'd3542,-16'd2248,16'd2883,16'd3817,16'd637,16'd3967,16'd1814,-16'd8336,-16'd6868,16'd3355,-16'd515,16'd3087,-16'd21,16'd1424,16'd1404};
dout[617]={ 16'd2096,-16'd958,16'd4315,-16'd5159,-16'd379,16'd6174,-16'd837,-16'd3064,-16'd3614,-16'd5533,-16'd814,-16'd660,-16'd742,-16'd153,-16'd1161,-16'd3528,16'd1020,-16'd295,-16'd2910,-16'd9873,-16'd3843,16'd3228,16'd368,16'd6231,-16'd919,16'd2324,16'd3082,16'd3082,16'd1651,16'd6219,-16'd5174,16'd2591,-16'd3786,-16'd4154,-16'd1777,-16'd4194};
dout[618]={ -16'd1533,-16'd6035,-16'd5280,-16'd6631,-16'd2817,-16'd5066,16'd558,16'd6313,-16'd3330,16'd1706,16'd3662,-16'd3215,-16'd4247,16'd1844,-16'd2616,-16'd6914,-16'd3743,-16'd2535,-16'd3928,16'd3810,-16'd3241,-16'd1788,16'd5134,-16'd4843,-16'd5770,-16'd2168,16'd1518,16'd614,-16'd3917,-16'd946,16'd6884,16'd2237,-16'd1550,-16'd3582,-16'd4606,-16'd3009};
dout[619]={ -16'd6253,-16'd874,16'd6150,16'd4242,16'd6259,16'd2071,-16'd2711,-16'd4372,-16'd3492,-16'd252,-16'd3245,16'd5393,16'd2846,16'd2222,-16'd3640,-16'd2263,16'd5024,16'd3402,16'd940,16'd4333,16'd3306,-16'd7503,-16'd3292,-16'd1361,-16'd5178,-16'd3039,16'd6241,16'd5660,16'd5087,-16'd2830,16'd3900,-16'd154,-16'd1101,16'd405,16'd7125,-16'd5720};
dout[620]={ 16'd75,-16'd2958,-16'd7486,-16'd590,16'd2805,16'd2954,-16'd6728,-16'd833,-16'd987,16'd5031,16'd942,16'd9362,-16'd4281,16'd8558,16'd2819,-16'd867,-16'd6774,-16'd398,16'd5438,16'd3225,16'd3982,-16'd4058,16'd7333,-16'd9025,-16'd5707,-16'd927,16'd1040,-16'd2906,-16'd7417,16'd3106,-16'd9729,16'd4681,-16'd5474,16'd1419,-16'd6656,16'd3163};
dout[621]={ -16'd1771,16'd3514,16'd2074,-16'd5772,16'd1171,16'd6012,-16'd1487,-16'd2641,16'd6012,16'd5594,16'd2839,-16'd2785,-16'd5489,16'd3357,16'd6159,16'd1681,-16'd792,-16'd3094,-16'd232,-16'd4684,-16'd1004,16'd3632,-16'd7053,-16'd7968,-16'd6761,16'd4836,16'd7564,16'd8236,-16'd1443,16'd6816,16'd3344,-16'd1540,16'd563,16'd2043,-16'd927,-16'd7067};
dout[622]={ 16'd8415,16'd7287,16'd3075,-16'd7678,16'd6095,-16'd1193,16'd3309,16'd6603,-16'd6326,-16'd2742,16'd1232,-16'd6291,16'd6895,-16'd3632,-16'd3204,16'd8800,-16'd1347,-16'd1463,16'd5690,16'd2477,16'd4040,-16'd3441,-16'd8194,16'd1281,-16'd7199,-16'd8918,16'd953,16'd2202,16'd3865,16'd3583,16'd4642,-16'd566,-16'd8316,-16'd1831,16'd6149,16'd3708};
dout[623]={ 16'd135,-16'd701,16'd1493,16'd633,16'd720,-16'd8353,-16'd6946,-16'd3426,-16'd7543,-16'd2425,-16'd13913,-16'd3588,-16'd6430,-16'd1479,-16'd3222,-16'd4511,16'd4127,-16'd7588,16'd2105,-16'd6092,16'd6768,-16'd11203,-16'd5982,16'd1410,-16'd3605,-16'd714,16'd4415,16'd7918,-16'd5811,-16'd702,16'd2533,-16'd4349,16'd2557,16'd544,-16'd3081,16'd1376};
dout[624]={ -16'd4340,-16'd4382,-16'd4151,-16'd7683,16'd3358,-16'd2797,-16'd453,-16'd63,-16'd270,16'd2064,-16'd7979,-16'd1406,-16'd4518,-16'd7529,16'd2188,-16'd8754,-16'd6813,-16'd8186,16'd5416,16'd5361,-16'd5771,-16'd2330,16'd4713,-16'd941,16'd4034,-16'd3263,-16'd8045,16'd533,-16'd8620,16'd4341,16'd6261,16'd8644,-16'd8544,-16'd6764,-16'd6808,-16'd5421};
dout[625]={ -16'd3403,16'd3472,-16'd2013,16'd921,-16'd4658,16'd5388,-16'd2032,16'd4777,16'd4591,-16'd3241,-16'd3860,-16'd1152,-16'd3010,-16'd2832,16'd4709,-16'd4098,16'd1701,16'd682,-16'd3382,-16'd3200,-16'd3767,-16'd6703,-16'd4116,16'd726,-16'd3098,-16'd554,-16'd5898,16'd6323,16'd1441,16'd4299,16'd2159,-16'd4338,-16'd4030,16'd4190,-16'd1541,16'd516};
dout[626]={ -16'd2874,16'd1839,16'd767,-16'd5535,-16'd2155,16'd6183,16'd5546,16'd2968,16'd5251,-16'd2966,-16'd637,16'd277,-16'd3236,16'd1595,16'd1513,16'd4371,-16'd1724,16'd3351,16'd2049,16'd62,-16'd55,-16'd3665,16'd413,-16'd3642,-16'd2304,16'd423,16'd275,16'd4871,16'd5820,-16'd1867,-16'd1364,-16'd3928,-16'd8744,-16'd6637,-16'd3025,16'd6379};
dout[627]={ 16'd272,16'd4533,16'd3362,-16'd1189,16'd2244,16'd4046,-16'd3826,-16'd1142,-16'd3150,16'd5210,-16'd680,-16'd6241,-16'd5000,-16'd1263,-16'd990,16'd2360,-16'd161,16'd6845,16'd3944,-16'd6447,-16'd1249,-16'd6239,16'd2381,16'd4229,-16'd6192,16'd478,16'd6078,-16'd5558,-16'd7641,16'd3807,16'd6197,-16'd5588,-16'd987,16'd2793,-16'd1140,-16'd2421};
dout[628]={ -16'd1328,16'd3231,16'd2260,-16'd853,-16'd4841,-16'd5939,-16'd4411,16'd538,-16'd3768,-16'd916,-16'd6689,-16'd5598,-16'd4959,16'd4024,-16'd275,-16'd6945,-16'd7514,-16'd1833,-16'd2878,-16'd6057,16'd3842,16'd1177,16'd3317,16'd5468,-16'd5052,16'd6415,-16'd852,-16'd5946,16'd883,16'd1855,-16'd4820,-16'd6207,-16'd2390,16'd1291,-16'd4011,-16'd4455};
dout[629]={ 16'd642,16'd3100,-16'd1805,16'd5339,16'd4632,16'd6281,16'd5894,16'd4225,-16'd762,16'd682,-16'd4532,-16'd5123,16'd4134,16'd3136,-16'd2605,16'd114,16'd4780,-16'd4117,16'd3776,16'd1183,-16'd2051,-16'd7524,16'd5464,16'd5733,-16'd6464,16'd3255,-16'd3149,-16'd3599,-16'd5975,16'd2507,16'd4289,-16'd4442,-16'd4703,16'd4726,16'd5475,-16'd4421};
dout[630]={ 16'd7002,16'd7828,16'd2397,-16'd2703,-16'd6748,16'd1361,16'd4727,16'd167,16'd8423,-16'd2295,16'd1117,-16'd2604,-16'd1266,-16'd4751,-16'd490,-16'd4206,-16'd2819,-16'd106,-16'd6008,16'd1284,16'd4318,16'd3183,16'd1218,-16'd8224,-16'd4425,-16'd11682,16'd2483,16'd8164,16'd6717,16'd2372,-16'd7391,16'd3948,16'd898,-16'd3331,-16'd11543,-16'd4494};
dout[631]={ 16'd417,-16'd7167,16'd2353,16'd1412,16'd5344,-16'd8040,-16'd6220,16'd1385,16'd8483,-16'd3969,-16'd500,16'd7222,-16'd7972,16'd4237,16'd8091,-16'd400,16'd5375,16'd6779,16'd4387,16'd96,16'd5714,16'd340,16'd6412,-16'd2988,-16'd5605,16'd4717,-16'd4480,16'd8479,-16'd2131,-16'd4082,-16'd5942,-16'd4088,-16'd9607,-16'd8227,16'd6997,-16'd126};
dout[632]={ 16'd2146,16'd2758,-16'd5206,16'd1103,16'd985,16'd145,16'd6358,-16'd6360,-16'd1667,-16'd6603,-16'd7319,-16'd6002,-16'd811,-16'd5259,-16'd289,16'd8649,16'd1053,-16'd1153,16'd6552,16'd3115,-16'd2643,16'd4202,-16'd6111,-16'd6798,-16'd5686,-16'd2844,-16'd5528,-16'd4577,16'd6023,-16'd2058,16'd1185,-16'd2073,-16'd7792,-16'd6162,16'd6675,-16'd7979};
dout[633]={ 16'd4544,16'd3615,-16'd2047,-16'd8203,-16'd6520,-16'd5495,-16'd7368,-16'd3717,16'd7024,16'd1762,-16'd13648,16'd7180,-16'd3349,-16'd1444,16'd1268,-16'd4160,16'd423,-16'd3567,16'd5843,-16'd807,-16'd5162,-16'd100,16'd6914,16'd4694,-16'd6128,-16'd782,16'd3396,16'd2313,-16'd1154,-16'd1571,-16'd7029,16'd3352,16'd1534,16'd1305,16'd37,-16'd7148};
dout[634]={ -16'd6841,16'd3733,16'd6968,-16'd2954,16'd381,-16'd2641,-16'd4932,-16'd2495,-16'd4721,-16'd8019,-16'd5395,16'd7692,16'd1542,-16'd1356,-16'd1049,16'd2867,16'd569,-16'd5311,-16'd6470,-16'd3002,16'd2982,-16'd9203,-16'd5968,-16'd829,-16'd4020,-16'd7338,16'd4179,-16'd1688,-16'd3869,16'd469,16'd1740,16'd103,16'd3876,-16'd2957,-16'd5782,16'd3885};
dout[635]={ -16'd4363,16'd6480,-16'd6317,16'd638,-16'd4263,-16'd6095,16'd6583,16'd3227,-16'd1022,-16'd3609,-16'd1778,16'd6409,16'd3435,-16'd3511,-16'd1659,-16'd6616,16'd1116,-16'd2925,16'd6195,-16'd6242,-16'd4526,-16'd4062,-16'd803,-16'd193,16'd473,-16'd3757,16'd2623,-16'd1289,16'd860,-16'd6955,-16'd1669,16'd7726,16'd2941,-16'd8482,16'd5463,16'd7247};
dout[636]={ 16'd1923,16'd2659,16'd5713,16'd6399,-16'd5799,-16'd6869,-16'd3815,-16'd1601,16'd603,16'd1120,16'd3417,-16'd2685,-16'd4148,-16'd2332,-16'd4478,-16'd4255,-16'd392,-16'd1037,16'd905,-16'd4716,-16'd5602,-16'd1166,-16'd4865,-16'd1516,16'd5334,-16'd31,-16'd8321,-16'd1992,-16'd4079,16'd1990,-16'd1136,-16'd4983,16'd4059,16'd595,16'd3634,16'd4302};
dout[637]={ -16'd4406,-16'd2821,-16'd8029,-16'd1082,16'd2511,16'd524,-16'd4519,16'd7748,-16'd6949,-16'd4489,-16'd5408,16'd5735,16'd4332,-16'd4077,-16'd4240,16'd5915,16'd4825,-16'd802,16'd6723,16'd415,16'd7050,-16'd3687,-16'd2798,16'd456,-16'd7021,16'd7256,-16'd1027,16'd928,-16'd7849,-16'd1482,-16'd1932,16'd5806,-16'd1417,16'd2198,-16'd5090,-16'd1340};
dout[638]={ 16'd3014,16'd6221,-16'd672,16'd5682,-16'd3094,16'd6869,-16'd1553,16'd5937,-16'd5775,16'd1075,16'd5804,16'd2553,16'd8809,16'd5254,16'd2226,-16'd4310,-16'd4108,16'd2531,16'd6807,-16'd2602,16'd682,16'd346,-16'd8259,16'd1461,-16'd7176,16'd4529,-16'd3016,16'd1307,16'd3400,-16'd1358,-16'd7068,-16'd6135,16'd606,-16'd1147,-16'd1760,16'd4838};
dout[639]={ 16'd22,16'd3023,16'd4831,-16'd3072,16'd4987,16'd1496,16'd1913,-16'd769,16'd1988,-16'd2862,16'd5880,-16'd166,-16'd2633,16'd1113,16'd3440,16'd5063,16'd3672,16'd5900,16'd1050,16'd753,16'd2394,16'd5774,-16'd1550,-16'd1952,-16'd7696,-16'd5207,16'd813,16'd582,16'd1649,16'd4948,16'd4699,16'd2670,-16'd3970,-16'd721,-16'd659,16'd6922};
dout[640]={ 16'd4333,16'd9793,-16'd2737,-16'd4011,-16'd8185,-16'd7080,-16'd5537,-16'd6998,16'd9603,-16'd4171,-16'd842,16'd2762,-16'd1304,-16'd2896,16'd3272,-16'd7977,16'd5226,-16'd4872,-16'd3277,16'd5253,16'd7402,-16'd1972,-16'd7208,-16'd5793,16'd2143,-16'd4702,16'd2573,16'd245,-16'd3620,16'd5676,-16'd7398,-16'd400,-16'd376,-16'd2040,-16'd2496,16'd6200};
dout[641]={ -16'd4665,-16'd1263,16'd3982,16'd542,-16'd5788,-16'd6162,-16'd6272,16'd5429,16'd6549,-16'd7438,16'd1811,16'd6366,-16'd6285,16'd6650,-16'd6852,16'd4129,-16'd4417,16'd5623,16'd2751,-16'd8531,16'd3197,16'd7443,16'd3653,16'd1853,-16'd2089,-16'd40,16'd5234,16'd4835,-16'd3611,-16'd978,-16'd226,-16'd3134,16'd1223,16'd5259,-16'd2534,-16'd6262};
dout[642]={ 16'd449,16'd3724,-16'd2038,16'd1366,-16'd3343,16'd1651,-16'd1801,16'd6211,-16'd597,16'd4181,-16'd2948,-16'd821,16'd3466,16'd8406,-16'd6155,16'd5637,16'd2781,16'd4626,-16'd1179,-16'd740,-16'd2669,16'd6055,-16'd7633,-16'd10284,16'd5033,-16'd5773,-16'd2906,16'd3027,-16'd3450,16'd7201,16'd3698,16'd1658,-16'd2801,-16'd5514,16'd10650,16'd5845};
dout[643]={ -16'd1606,16'd988,-16'd7341,16'd1353,-16'd6817,-16'd1273,16'd3655,16'd5712,16'd51,-16'd3976,-16'd2426,16'd8983,16'd1527,-16'd5102,16'd6584,16'd2596,16'd2635,-16'd8831,16'd7712,16'd207,16'd6139,-16'd5922,-16'd4274,16'd392,16'd1267,-16'd9158,-16'd8644,-16'd864,16'd3580,-16'd199,16'd3882,-16'd2391,16'd2317,-16'd5635,-16'd365,-16'd6892};
dout[644]={ 16'd6498,-16'd5552,-16'd2084,-16'd4481,-16'd4661,16'd1599,-16'd5632,16'd3174,16'd1093,-16'd3217,-16'd11503,-16'd1831,16'd5193,16'd3465,-16'd1319,16'd5124,16'd18,-16'd7468,-16'd6299,-16'd7281,-16'd4049,-16'd3996,-16'd1476,-16'd69,-16'd4656,-16'd6181,-16'd1157,16'd7517,-16'd9580,-16'd3678,-16'd3545,16'd6046,-16'd3895,16'd2674,-16'd8586,-16'd5246};
dout[645]={ 16'd2433,16'd3598,-16'd2024,-16'd8033,16'd3521,16'd3790,16'd4360,16'd3065,-16'd1714,16'd1917,16'd3061,-16'd1546,16'd3482,16'd5276,-16'd2488,-16'd8303,-16'd4465,-16'd1538,-16'd2372,16'd8763,-16'd5382,16'd4526,16'd5225,-16'd5421,16'd4128,-16'd1950,-16'd919,16'd1948,16'd3861,-16'd2445,16'd1619,16'd1038,16'd808,-16'd4873,-16'd6268,16'd5897};
dout[646]={ 16'd122,-16'd5553,16'd5638,-16'd6183,-16'd2215,16'd4714,-16'd3373,-16'd6438,16'd4692,16'd3683,-16'd5884,-16'd3128,16'd2417,-16'd3071,16'd3197,-16'd5992,16'd5192,16'd5137,16'd1445,-16'd1950,16'd3863,-16'd2029,-16'd4782,-16'd2588,16'd1684,16'd5631,16'd5653,16'd3,-16'd7667,-16'd2005,16'd2200,-16'd634,16'd4438,-16'd2437,16'd2873,-16'd6994};
dout[647]={ -16'd6868,-16'd5243,-16'd537,-16'd5575,16'd4805,16'd3029,-16'd227,-16'd1247,-16'd4653,-16'd151,16'd4408,-16'd1253,16'd7540,-16'd3839,-16'd816,16'd7311,16'd3493,-16'd7505,16'd6166,16'd348,-16'd1387,16'd373,-16'd5528,16'd1351,16'd4290,16'd5061,16'd3703,16'd989,16'd5123,-16'd1107,-16'd2954,-16'd2224,-16'd1336,-16'd1949,16'd2144,16'd7658};
dout[648]={ 16'd5457,16'd5864,16'd6063,16'd1555,-16'd651,-16'd6646,16'd864,-16'd5568,16'd2122,16'd271,-16'd3210,-16'd4756,16'd6761,-16'd4989,-16'd3699,-16'd4537,-16'd1963,-16'd2369,16'd5306,-16'd4219,16'd4619,-16'd8590,-16'd3481,-16'd1674,16'd6444,16'd1873,-16'd8269,16'd6258,16'd5514,-16'd348,16'd3054,16'd444,-16'd3245,16'd2609,-16'd1956,-16'd1149};
dout[649]={ 16'd2615,16'd1899,16'd623,-16'd6988,16'd1810,-16'd2643,16'd821,-16'd4755,16'd161,-16'd3854,16'd5651,16'd675,-16'd4914,16'd1069,16'd7415,-16'd5772,-16'd912,16'd1415,16'd7693,-16'd6765,-16'd95,-16'd6292,16'd6091,16'd5684,-16'd5811,-16'd4231,16'd3094,-16'd1705,16'd438,16'd2432,16'd886,16'd6832,16'd2811,-16'd3767,16'd5864,-16'd5744};
dout[650]={ -16'd7069,16'd6385,-16'd4298,16'd2084,-16'd10980,16'd1423,-16'd7332,-16'd1721,-16'd706,-16'd1700,16'd4553,-16'd6028,16'd4653,-16'd1560,-16'd7094,-16'd1836,16'd2731,16'd2494,16'd2741,16'd6324,-16'd3023,-16'd3620,-16'd8696,16'd2844,16'd2810,16'd3307,-16'd3075,16'd337,16'd4639,-16'd5360,16'd2894,-16'd8874,-16'd5761,-16'd3556,16'd1550,-16'd8232};
dout[651]={ -16'd4872,-16'd2658,16'd4062,-16'd4906,-16'd5125,-16'd5434,-16'd3859,-16'd4073,16'd2184,16'd7732,-16'd52,16'd5694,-16'd8984,16'd997,-16'd5434,16'd1787,16'd1476,16'd2916,-16'd5103,16'd790,16'd1719,16'd3210,-16'd4387,-16'd5358,-16'd6679,16'd9301,-16'd2317,16'd2565,16'd4147,-16'd8061,16'd943,16'd4341,-16'd2414,16'd6696,16'd7704,-16'd2524};
dout[652]={ -16'd7748,-16'd4092,16'd1966,16'd2225,-16'd7274,16'd5321,16'd913,-16'd9866,16'd1690,16'd1647,16'd1050,16'd4144,16'd4902,-16'd953,16'd746,-16'd2554,-16'd7892,-16'd561,16'd611,16'd1758,-16'd4953,16'd4540,16'd5867,-16'd6235,16'd2773,-16'd655,-16'd141,16'd9438,16'd4184,-16'd2042,16'd1868,16'd146,-16'd3874,16'd5932,16'd9159,-16'd1135};
dout[653]={ 16'd1321,-16'd11342,16'd3813,16'd140,16'd1526,-16'd5784,-16'd4810,-16'd4041,-16'd1240,-16'd5050,-16'd7728,16'd5269,16'd3919,16'd5084,-16'd6058,16'd5949,-16'd5101,-16'd6799,-16'd5489,16'd1476,16'd3304,-16'd7165,16'd203,16'd3512,-16'd9793,-16'd12586,-16'd4195,16'd7559,16'd7987,16'd1272,-16'd8244,16'd1098,-16'd8033,-16'd5915,16'd2067,-16'd4483};
dout[654]={ 16'd1743,-16'd5026,-16'd5307,-16'd8750,-16'd1600,16'd2519,16'd5742,-16'd3843,16'd1645,-16'd1183,-16'd9851,-16'd2310,-16'd5951,-16'd3900,16'd1112,16'd6360,-16'd8550,-16'd2914,16'd548,-16'd2751,-16'd4343,-16'd5628,-16'd2223,16'd2491,-16'd7638,-16'd3614,-16'd4241,16'd1234,-16'd665,16'd3074,-16'd6620,16'd4092,-16'd6421,16'd3901,16'd456,-16'd7652};
dout[655]={ -16'd7647,16'd6875,-16'd5346,16'd5257,16'd2403,-16'd8058,16'd4517,-16'd1744,-16'd950,16'd871,-16'd8861,16'd4078,-16'd4738,-16'd406,16'd4662,16'd3198,-16'd6651,16'd1450,16'd2426,-16'd755,16'd1695,-16'd6217,16'd5263,16'd2201,-16'd389,16'd5142,-16'd1754,-16'd5244,16'd2186,-16'd3448,16'd213,-16'd636,-16'd3074,16'd4380,16'd4437,-16'd7147};
dout[656]={ -16'd4462,16'd7322,-16'd2810,-16'd7761,16'd2526,-16'd102,-16'd818,-16'd5849,16'd4831,16'd1525,16'd883,16'd527,-16'd6405,16'd6693,-16'd4070,-16'd1660,-16'd2743,-16'd5884,16'd7356,-16'd3559,-16'd3960,16'd6256,-16'd5182,16'd1855,-16'd5308,-16'd167,-16'd5765,-16'd2137,-16'd5068,-16'd3261,-16'd4394,-16'd2288,-16'd381,-16'd1000,16'd492,16'd2761};
dout[657]={ 16'd2500,16'd6942,-16'd590,16'd5570,16'd6352,-16'd860,-16'd4924,16'd715,-16'd4769,16'd856,-16'd1768,-16'd7550,-16'd51,16'd6344,16'd4050,-16'd4440,16'd1560,-16'd4919,-16'd4549,16'd3656,-16'd4098,16'd2008,-16'd834,16'd5200,-16'd1513,-16'd5207,16'd2479,-16'd1330,16'd1391,16'd4218,-16'd1583,16'd3070,-16'd982,-16'd5449,16'd279,-16'd5668};
dout[658]={ 16'd702,-16'd7994,16'd692,-16'd2105,16'd6983,16'd1422,-16'd5380,-16'd2054,-16'd5047,16'd2535,16'd1666,16'd5802,-16'd4535,16'd5000,-16'd1200,16'd6155,-16'd3937,-16'd4888,16'd10594,-16'd3304,-16'd3069,16'd1609,-16'd6944,-16'd580,-16'd4928,16'd2480,16'd5592,16'd6568,-16'd8850,16'd6006,16'd6647,-16'd687,-16'd5587,16'd203,-16'd1783,16'd5452};
dout[659]={ -16'd7583,-16'd5580,16'd2188,16'd6634,16'd4513,-16'd3397,16'd1114,16'd4944,16'd373,16'd1433,-16'd6733,-16'd3854,16'd6328,-16'd220,16'd427,-16'd699,-16'd1645,-16'd5106,-16'd2772,16'd2492,16'd5100,-16'd4286,-16'd1648,16'd3498,16'd355,-16'd4702,16'd3920,-16'd5534,-16'd1880,16'd12,16'd476,-16'd4332,16'd247,16'd998,-16'd1391,-16'd2036};
dout[660]={ -16'd3129,-16'd1675,-16'd1271,-16'd1677,-16'd8632,-16'd7174,-16'd2454,16'd622,16'd1961,16'd1325,16'd3743,-16'd5275,16'd8382,-16'd5344,16'd1415,16'd5799,-16'd6057,-16'd57,16'd474,-16'd1060,-16'd12071,16'd9307,-16'd2899,16'd2258,16'd4260,-16'd3787,16'd1990,-16'd3816,-16'd4134,-16'd5854,-16'd5856,16'd1789,-16'd1936,-16'd3757,-16'd7546,16'd1321};
dout[661]={ 16'd819,-16'd5065,-16'd337,-16'd8868,16'd2624,-16'd1700,16'd1995,-16'd4131,16'd8351,16'd7743,16'd7938,16'd5389,-16'd371,16'd5370,-16'd5946,-16'd6516,-16'd4193,16'd3888,16'd2291,16'd2681,-16'd1537,16'd6455,-16'd1796,-16'd6654,-16'd5145,16'd2579,-16'd1311,16'd7003,16'd3685,-16'd2721,-16'd1228,16'd3771,-16'd3769,-16'd5330,-16'd208,-16'd7964};
dout[662]={ -16'd1880,-16'd1258,-16'd2219,-16'd7877,16'd203,-16'd7996,-16'd5167,-16'd6649,16'd6552,16'd5018,-16'd662,16'd1093,-16'd788,16'd6977,16'd2005,16'd5505,16'd724,-16'd318,-16'd4534,16'd5285,16'd2245,-16'd1727,-16'd7948,-16'd761,16'd4302,16'd5702,-16'd4236,16'd5520,-16'd4159,-16'd7091,16'd3746,16'd8094,16'd6271,-16'd8728,16'd4717,16'd4331};
dout[663]={ 16'd668,-16'd2147,16'd5265,-16'd8069,-16'd233,16'd6434,16'd2398,16'd3741,-16'd8632,-16'd3535,-16'd6178,-16'd6228,-16'd25,16'd8728,16'd5199,-16'd4480,16'd4039,-16'd1628,16'd263,16'd7919,-16'd2738,16'd1015,16'd4614,16'd1506,16'd5131,-16'd15229,-16'd1797,16'd8506,-16'd1833,16'd5519,-16'd1195,16'd681,16'd6072,16'd610,16'd2258,-16'd4698};
dout[664]={ -16'd154,16'd951,-16'd138,-16'd3340,-16'd4423,-16'd286,-16'd1304,-16'd642,16'd891,-16'd5519,-16'd4736,16'd1083,-16'd4409,-16'd299,-16'd4815,16'd4679,16'd5745,16'd733,-16'd5212,16'd838,-16'd504,16'd3804,16'd1883,16'd5093,16'd4683,-16'd3986,16'd1458,16'd5778,-16'd3442,16'd173,16'd1071,-16'd5855,-16'd2237,-16'd5582,-16'd45,-16'd920};
dout[665]={ 16'd5713,-16'd4216,-16'd3700,-16'd6085,16'd5523,16'd4221,-16'd4698,16'd1625,-16'd37,16'd5171,-16'd223,-16'd5475,-16'd8363,16'd3952,-16'd3795,-16'd500,-16'd3778,16'd369,16'd106,-16'd3884,16'd1403,-16'd4552,-16'd8452,16'd3192,-16'd1578,16'd6717,-16'd249,16'd148,16'd4061,16'd724,16'd3947,16'd1150,-16'd5369,16'd3966,-16'd2401,16'd6771};
dout[666]={ -16'd1044,-16'd4544,16'd4205,16'd5620,16'd1368,-16'd482,-16'd1910,16'd124,-16'd42,-16'd742,16'd1011,-16'd523,-16'd4391,16'd1505,-16'd481,-16'd4688,16'd6504,16'd1946,-16'd5621,16'd3091,16'd1362,-16'd4197,-16'd2980,-16'd3485,16'd5621,16'd2410,-16'd1604,16'd4871,-16'd519,-16'd5810,-16'd5107,16'd379,16'd6598,-16'd235,-16'd3240,-16'd2232};
dout[667]={ -16'd1784,-16'd998,16'd2816,16'd756,-16'd5843,16'd1279,16'd1968,-16'd6366,16'd7194,16'd471,16'd1201,-16'd5111,-16'd6497,-16'd5747,16'd7119,-16'd3383,-16'd3899,16'd1662,16'd6592,16'd4053,16'd1302,-16'd3870,-16'd1735,16'd4394,-16'd3719,-16'd3641,-16'd5913,16'd1543,16'd4205,16'd6831,-16'd2489,16'd3749,16'd56,-16'd5892,16'd6523,16'd32};
dout[668]={ 16'd5363,-16'd6299,16'd5989,-16'd2908,16'd5169,16'd3365,16'd3829,-16'd2918,-16'd2340,16'd5260,-16'd3032,-16'd1692,16'd1770,-16'd6322,16'd6872,16'd7087,16'd5294,-16'd6078,16'd5345,-16'd2191,16'd3266,16'd1687,-16'd3498,-16'd3990,-16'd6378,-16'd3509,-16'd4572,-16'd3740,16'd2882,16'd2012,16'd2573,16'd1936,16'd6085,-16'd2020,-16'd3856,-16'd3532};
dout[669]={ -16'd7884,16'd5588,16'd2,16'd5552,16'd2236,-16'd5745,16'd2276,16'd7592,16'd4076,16'd1406,-16'd3017,16'd3883,16'd5780,16'd1741,-16'd2885,-16'd2223,16'd331,16'd2698,16'd2458,16'd2180,-16'd6378,16'd4703,-16'd1560,16'd5644,-16'd8810,16'd5460,-16'd5866,16'd6828,-16'd3328,16'd2056,-16'd5248,16'd4221,-16'd5218,16'd456,-16'd1237,16'd3907};
dout[670]={ 16'd2436,16'd7986,-16'd2637,-16'd2828,16'd3674,-16'd105,-16'd1121,-16'd378,16'd10087,16'd605,16'd4895,-16'd2385,16'd3104,16'd9798,-16'd2834,-16'd1528,16'd4372,-16'd3885,16'd4332,-16'd1536,-16'd12952,16'd1670,16'd1864,16'd7611,16'd3458,16'd1646,-16'd1161,16'd6123,-16'd3680,16'd216,-16'd5827,16'd1174,-16'd8133,-16'd4409,-16'd1457,-16'd9175};
dout[671]={ -16'd9174,16'd382,-16'd6597,16'd5013,16'd6428,-16'd502,-16'd2353,-16'd3360,16'd976,16'd5339,16'd2434,16'd3726,16'd1165,16'd5504,16'd2749,-16'd4042,16'd1009,-16'd6284,16'd2536,16'd9281,-16'd4273,16'd11738,-16'd6665,-16'd3484,-16'd6693,16'd10503,-16'd2558,16'd396,16'd6055,-16'd4836,-16'd43,16'd411,-16'd5176,16'd5504,-16'd2493,-16'd8225};
dout[672]={ 16'd6171,-16'd5213,-16'd2443,-16'd5583,-16'd5970,16'd2495,-16'd78,16'd4517,16'd410,16'd1624,-16'd6268,16'd9222,16'd3502,16'd8107,-16'd1360,-16'd5123,16'd3289,16'd3506,16'd2314,-16'd2183,-16'd3292,16'd787,16'd3836,-16'd1529,16'd4592,-16'd1045,16'd6076,16'd4810,-16'd6352,-16'd650,16'd3890,16'd580,-16'd7215,16'd4132,16'd1224,16'd1946};
dout[673]={ 16'd1203,16'd1377,-16'd7443,-16'd96,-16'd780,16'd3498,16'd323,16'd3819,-16'd7128,-16'd4388,16'd2154,-16'd7026,16'd2061,16'd11715,-16'd5834,16'd7015,-16'd7676,-16'd2286,-16'd3175,16'd6019,16'd1441,-16'd5312,16'd1194,16'd632,-16'd4811,-16'd13404,16'd4503,16'd10112,16'd8684,-16'd5036,-16'd3878,16'd3582,-16'd3377,-16'd476,16'd8020,16'd5614};
dout[674]={ 16'd3075,-16'd804,-16'd2610,-16'd6428,-16'd1935,-16'd3732,16'd6912,-16'd2444,16'd4361,16'd4858,16'd5974,-16'd7997,-16'd4826,16'd6788,-16'd2984,16'd8170,-16'd7105,16'd6537,-16'd4321,16'd7612,16'd2794,16'd1522,16'd4931,-16'd5840,16'd6283,-16'd5036,16'd4878,-16'd1851,16'd4237,16'd4502,-16'd6262,-16'd1217,16'd831,16'd6580,-16'd3408,16'd5955};
dout[675]={ -16'd3775,-16'd5326,-16'd5986,16'd3033,16'd1262,-16'd4679,16'd1731,-16'd3636,-16'd3579,16'd2842,-16'd4608,-16'd3938,-16'd6101,16'd5724,-16'd5880,16'd1567,-16'd5628,-16'd2150,16'd3045,16'd3427,-16'd4770,16'd3851,16'd5979,-16'd21,-16'd6947,-16'd1887,-16'd5770,-16'd927,16'd6,16'd2122,16'd1218,-16'd202,-16'd5454,-16'd4852,-16'd6192,16'd226};
dout[676]={ 16'd399,-16'd1167,-16'd90,16'd4324,-16'd6803,16'd2227,16'd3916,-16'd5781,-16'd3585,16'd1463,16'd2423,16'd4171,16'd369,-16'd5170,16'd5814,16'd2566,16'd543,-16'd4493,-16'd4791,16'd712,-16'd3976,16'd4439,-16'd6550,16'd5397,16'd567,16'd371,-16'd2841,16'd4088,16'd659,16'd7406,16'd2100,-16'd5111,-16'd6077,-16'd3854,-16'd808,16'd3632};
dout[677]={ -16'd3284,-16'd4137,16'd5501,-16'd6955,-16'd5747,-16'd3212,-16'd4484,-16'd2668,16'd5895,16'd4098,16'd4684,16'd3054,16'd424,-16'd411,16'd4349,16'd762,-16'd2396,-16'd7534,16'd1457,16'd1438,-16'd3387,16'd4650,16'd5382,-16'd449,-16'd5140,16'd5560,16'd5804,-16'd3766,-16'd7563,-16'd2569,-16'd6521,16'd1098,-16'd5102,16'd50,16'd8723,16'd7053};
dout[678]={ -16'd8371,-16'd4700,-16'd3215,-16'd1271,-16'd1194,16'd2062,-16'd3941,16'd7202,16'd676,16'd924,16'd3339,-16'd8373,-16'd2934,-16'd3895,-16'd2215,-16'd5173,16'd2006,-16'd164,-16'd2198,-16'd2865,16'd1578,-16'd6889,-16'd8836,16'd7968,16'd6435,-16'd4920,16'd5356,-16'd4031,16'd5651,-16'd3070,16'd1174,16'd3185,16'd1748,-16'd6802,16'd3717,16'd2514};
dout[679]={ -16'd6210,16'd2670,-16'd7628,-16'd7308,-16'd2231,-16'd3416,-16'd3105,-16'd2417,-16'd6095,-16'd2528,16'd2218,16'd3502,-16'd6511,16'd5573,-16'd2591,16'd3244,16'd2358,16'd3862,16'd2413,-16'd5629,16'd2652,-16'd1463,-16'd3655,16'd2386,16'd5900,16'd3493,16'd3165,-16'd2543,-16'd4131,-16'd4118,-16'd5752,16'd4544,16'd6036,-16'd6058,16'd900,16'd1065};
dout[680]={ -16'd36,-16'd243,16'd3494,-16'd4044,16'd5582,-16'd2250,16'd8392,-16'd7140,-16'd177,-16'd501,16'd4782,-16'd5767,16'd5535,16'd4983,-16'd3102,-16'd3935,-16'd3369,-16'd8063,-16'd4542,-16'd8680,-16'd6062,16'd4397,16'd2146,-16'd602,16'd5138,16'd10373,-16'd3188,16'd3969,-16'd1175,-16'd3068,16'd5072,16'd8636,-16'd8495,-16'd4031,-16'd3839,-16'd6655};
dout[681]={ -16'd7721,-16'd6279,-16'd2943,16'd1303,16'd3930,-16'd8128,-16'd750,-16'd9378,16'd515,16'd2342,-16'd3362,16'd87,16'd5725,-16'd2557,16'd6145,-16'd7552,-16'd8435,16'd4387,16'd3643,-16'd1920,16'd3540,-16'd185,16'd812,16'd2106,-16'd790,16'd6196,-16'd4441,-16'd481,-16'd1971,-16'd4390,-16'd2386,-16'd2766,-16'd5053,16'd230,16'd29,16'd2842};
dout[682]={ -16'd1195,-16'd2725,-16'd9485,16'd5601,-16'd1100,-16'd4499,16'd3239,-16'd7505,16'd1519,-16'd7265,16'd334,-16'd3122,-16'd4163,16'd505,-16'd4654,-16'd2552,-16'd5965,16'd4439,16'd2880,-16'd5873,16'd6755,16'd4942,-16'd6567,-16'd5152,16'd4121,16'd4260,16'd5394,16'd7493,16'd3492,-16'd7439,16'd8517,-16'd417,-16'd7666,-16'd6555,16'd9253,16'd325};
dout[683]={ -16'd6801,-16'd9704,-16'd10589,-16'd1761,-16'd4793,-16'd5473,16'd4438,-16'd983,-16'd2145,-16'd8562,-16'd2153,16'd1324,-16'd544,16'd10958,-16'd3563,16'd4099,-16'd2532,16'd1562,-16'd1338,-16'd2717,16'd4516,16'd3837,-16'd5033,16'd4881,16'd6950,-16'd5893,-16'd4854,16'd10768,-16'd6193,-16'd4673,-16'd5216,-16'd3689,-16'd6120,16'd988,16'd4130,-16'd6735};
dout[684]={ 16'd862,-16'd3337,-16'd2008,-16'd1715,-16'd7974,-16'd8209,16'd3776,-16'd3466,16'd4736,-16'd7848,-16'd2676,16'd2066,16'd799,16'd1631,-16'd5918,-16'd272,-16'd2476,-16'd1682,16'd9497,16'd9678,-16'd5031,-16'd761,-16'd7160,-16'd6219,-16'd321,-16'd4244,-16'd5029,16'd7689,-16'd3357,-16'd1162,-16'd2679,16'd2810,-16'd8363,16'd6013,-16'd305,-16'd267};
dout[685]={ -16'd1594,-16'd6727,-16'd4017,-16'd6757,-16'd5592,16'd5052,-16'd980,16'd2262,-16'd1691,-16'd6953,16'd164,-16'd3271,-16'd9211,-16'd3481,16'd131,-16'd653,16'd1557,16'd6027,16'd3064,-16'd733,-16'd2655,-16'd3855,-16'd1467,-16'd1873,16'd830,16'd7619,16'd275,-16'd1363,-16'd3614,16'd8251,-16'd1645,-16'd1032,16'd1200,16'd1401,-16'd858,16'd3816};
dout[686]={ -16'd1524,-16'd4498,-16'd1902,-16'd6476,16'd5393,16'd70,16'd4774,-16'd5162,16'd4935,16'd2921,-16'd171,-16'd792,16'd4200,16'd5086,16'd295,-16'd2264,16'd6981,-16'd772,16'd42,16'd6131,16'd1677,-16'd1527,-16'd775,16'd1184,16'd1475,16'd1120,-16'd6587,-16'd3522,16'd3412,-16'd3645,16'd2508,-16'd2182,-16'd1468,-16'd5933,16'd5042,16'd2253};
dout[687]={ 16'd2820,-16'd3423,-16'd3514,-16'd4732,-16'd3013,-16'd2469,16'd6775,-16'd7560,-16'd5291,16'd315,16'd7412,16'd7557,-16'd7244,-16'd2955,-16'd7406,-16'd844,16'd8186,-16'd3363,16'd2278,-16'd492,-16'd3400,-16'd4006,-16'd7743,16'd1709,16'd4105,-16'd3672,-16'd3316,16'd8248,16'd6160,-16'd222,16'd4402,16'd3607,-16'd5860,-16'd2965,16'd1915,-16'd7280};
dout[688]={ -16'd1980,-16'd634,-16'd5284,-16'd5501,-16'd2472,-16'd4947,-16'd2913,-16'd6024,-16'd1087,16'd496,-16'd5996,-16'd6611,16'd1325,-16'd5834,16'd2483,-16'd4939,16'd4360,16'd5453,-16'd6025,-16'd512,16'd479,-16'd2101,-16'd2221,16'd3970,-16'd4193,16'd2271,-16'd6474,16'd190,16'd1827,16'd6642,-16'd8280,-16'd2116,-16'd4356,-16'd3767,16'd4281,-16'd5767};
dout[689]={ -16'd2439,-16'd2126,-16'd6758,16'd1911,-16'd6782,-16'd2917,16'd3001,-16'd6107,16'd1337,16'd1949,16'd2037,-16'd6074,-16'd69,-16'd762,-16'd6949,16'd4475,16'd3140,-16'd2145,-16'd3691,-16'd1879,-16'd2618,16'd5708,16'd3347,16'd7395,-16'd1038,16'd3541,-16'd1310,16'd7626,-16'd5311,16'd728,-16'd4852,16'd1100,-16'd7664,-16'd2764,-16'd3114,-16'd2926};
dout[690]={ -16'd3687,16'd3242,-16'd5250,16'd4925,16'd1871,-16'd9154,16'd4919,-16'd2625,16'd2863,-16'd802,16'd5441,-16'd4180,-16'd5235,16'd6234,16'd2663,16'd3342,-16'd6766,16'd4853,-16'd677,-16'd1889,16'd1115,-16'd191,16'd3025,16'd5971,-16'd274,16'd7403,-16'd3227,16'd8689,-16'd4521,16'd4645,16'd4670,16'd1677,16'd3081,16'd66,16'd4041,-16'd9203};
dout[691]={ -16'd5552,-16'd2309,16'd1763,16'd2688,16'd10354,16'd2736,16'd6326,-16'd5265,16'd8516,-16'd5793,-16'd1314,16'd4578,16'd6591,-16'd2059,16'd4701,-16'd4439,16'd5438,-16'd8369,16'd3485,16'd4668,16'd5194,16'd1579,-16'd5458,16'd166,16'd222,-16'd2697,16'd5343,16'd816,-16'd5394,16'd4043,16'd8123,-16'd487,-16'd5169,16'd4547,-16'd5566,-16'd5016};
dout[692]={ 16'd8064,16'd4964,16'd1504,16'd5564,16'd8304,16'd34,16'd6463,16'd5325,-16'd1028,-16'd7240,-16'd3508,-16'd2746,16'd381,16'd125,16'd10057,16'd7961,-16'd5467,16'd3460,16'd1563,16'd3153,16'd10672,16'd2857,-16'd1438,-16'd407,-16'd1378,-16'd981,16'd2865,16'd2410,16'd501,-16'd7555,16'd3418,-16'd4133,16'd5761,-16'd1850,16'd8355,16'd6596};
dout[693]={ -16'd7708,16'd5097,-16'd246,-16'd5018,-16'd2221,-16'd4139,16'd5357,16'd128,-16'd2335,-16'd9201,-16'd1059,-16'd9220,16'd1019,16'd300,-16'd2637,16'd3371,-16'd6188,16'd2560,16'd996,-16'd5065,16'd3176,16'd3193,-16'd667,16'd1027,-16'd5738,-16'd5839,-16'd988,-16'd2814,16'd5994,-16'd4212,16'd2790,16'd5706,16'd5314,-16'd1017,16'd3697,-16'd1847};
dout[694]={ -16'd8217,-16'd4144,-16'd8274,-16'd5921,16'd1898,-16'd8492,-16'd7447,-16'd4859,-16'd6424,16'd4937,16'd82,-16'd7548,-16'd3937,16'd7973,-16'd9431,16'd146,-16'd4491,-16'd2460,16'd3097,16'd6390,16'd3769,16'd3586,-16'd2084,16'd461,-16'd5137,16'd3602,-16'd4862,-16'd2306,16'd8059,16'd5646,-16'd5340,16'd5884,16'd380,16'd18,16'd253,-16'd4370};
dout[695]={ -16'd7143,-16'd7023,-16'd5534,-16'd323,16'd4219,-16'd4140,16'd1620,-16'd123,16'd7311,-16'd7563,16'd7836,-16'd5073,16'd2548,16'd3932,-16'd8619,16'd1823,-16'd8987,16'd6693,-16'd2129,-16'd3756,-16'd3218,-16'd1544,16'd2499,-16'd20,-16'd6014,-16'd5332,-16'd5795,16'd4347,-16'd7140,16'd2456,16'd1748,-16'd142,-16'd3871,-16'd6660,-16'd2496,-16'd2401};
dout[696]={ 16'd4870,-16'd8935,16'd9137,-16'd1147,-16'd1517,-16'd5907,-16'd6057,-16'd2374,-16'd1234,-16'd7043,-16'd2132,-16'd239,-16'd6026,16'd3176,-16'd5938,-16'd4057,-16'd4051,16'd5025,-16'd1067,-16'd7124,16'd5074,16'd2257,-16'd8162,16'd6635,16'd4861,-16'd5871,-16'd7741,16'd3345,16'd4598,-16'd4969,-16'd1696,16'd1623,16'd4037,16'd3843,16'd7523,16'd2287};
dout[697]={ 16'd4576,-16'd8302,16'd2327,16'd5070,16'd4213,16'd1188,16'd6822,16'd3208,-16'd135,-16'd4055,16'd3130,-16'd4424,-16'd5251,16'd4205,16'd4079,16'd5360,-16'd985,-16'd5702,-16'd7388,-16'd6243,-16'd4258,16'd4157,-16'd2981,-16'd909,-16'd5139,-16'd5498,-16'd7009,-16'd98,16'd3486,16'd5878,16'd2149,-16'd4227,-16'd799,-16'd4250,-16'd3900,-16'd7684};
dout[698]={ 16'd5859,16'd1427,-16'd2856,-16'd4667,16'd3386,-16'd7614,16'd5052,-16'd1071,16'd4225,16'd2395,16'd1063,-16'd704,16'd3978,-16'd6391,-16'd3373,-16'd5974,-16'd6604,16'd4924,16'd2793,16'd7475,16'd4697,16'd3567,16'd985,-16'd2939,-16'd914,-16'd6842,-16'd1297,-16'd3795,16'd7430,16'd542,-16'd4073,16'd3059,-16'd5302,-16'd2027,16'd2569,16'd6851};
dout[699]={ 16'd3442,-16'd3012,16'd3939,-16'd4256,-16'd7697,16'd7117,16'd1279,16'd3027,16'd6868,-16'd4725,-16'd163,16'd476,16'd4631,-16'd6049,16'd841,-16'd523,16'd933,-16'd6158,16'd1396,-16'd3687,16'd4470,-16'd4945,-16'd2144,-16'd5387,16'd1064,-16'd5687,16'd1421,-16'd1366,16'd3671,16'd1605,-16'd1871,-16'd3027,-16'd7467,16'd875,-16'd663,-16'd5447};
dout[700]={ 16'd3474,16'd1223,-16'd1209,-16'd5016,16'd4331,-16'd2518,16'd10545,-16'd2603,16'd6492,-16'd4139,16'd6009,-16'd1331,16'd5842,16'd5877,16'd4312,16'd10159,-16'd5265,16'd2102,-16'd1051,-16'd7845,16'd5992,16'd1538,-16'd3435,-16'd1209,-16'd8718,-16'd2606,-16'd2375,16'd9163,-16'd7892,-16'd700,-16'd911,16'd6872,-16'd5130,-16'd3718,-16'd8547,-16'd2357};
dout[701]={ -16'd1049,-16'd7618,-16'd11744,16'd4565,16'd5472,-16'd3483,-16'd565,-16'd2051,-16'd282,-16'd5582,16'd2021,16'd4716,-16'd2897,16'd1334,-16'd1545,16'd4168,16'd3609,-16'd837,16'd8104,-16'd3360,16'd7456,-16'd6749,16'd610,-16'd80,16'd4020,16'd3840,-16'd9220,-16'd4082,-16'd9111,16'd1642,-16'd356,-16'd4536,16'd1304,16'd4448,-16'd1701,16'd464};
dout[702]={ 16'd6825,16'd7322,-16'd10413,16'd6104,16'd5090,16'd6258,16'd7607,16'd5919,-16'd629,16'd2732,-16'd7714,-16'd1286,16'd9772,-16'd5616,-16'd3083,-16'd3622,16'd6150,-16'd9004,16'd8453,-16'd5723,16'd531,-16'd1639,16'd4361,16'd5989,-16'd7695,16'd7267,-16'd8144,-16'd4012,-16'd5270,-16'd5599,16'd2512,16'd2493,-16'd6407,16'd5201,16'd1678,-16'd1185};
dout[703]={ -16'd57,-16'd1829,-16'd13187,16'd4414,16'd5369,-16'd37,16'd2570,-16'd702,-16'd2412,-16'd1563,16'd2828,-16'd5629,16'd3629,16'd4264,16'd7488,16'd8976,-16'd4694,16'd858,16'd3161,16'd1633,-16'd954,-16'd1368,-16'd8524,16'd757,16'd65,-16'd3618,-16'd7994,-16'd1386,16'd359,16'd4220,16'd5571,16'd696,-16'd4231,-16'd5866,16'd3442,16'd5664};
dout[704]={ 16'd1496,-16'd2605,16'd864,16'd5765,-16'd5084,-16'd4350,16'd3599,-16'd8255,16'd5268,-16'd5603,16'd6116,16'd1741,16'd5171,16'd2938,16'd6011,16'd3292,-16'd7888,-16'd2989,-16'd1806,-16'd101,-16'd268,16'd7565,-16'd1355,16'd4146,-16'd1178,-16'd1535,-16'd1752,16'd356,16'd6966,16'd193,-16'd272,-16'd916,16'd505,-16'd1092,-16'd4834,16'd5503};
dout[705]={ -16'd1447,-16'd4069,16'd4284,-16'd4587,-16'd2104,16'd5003,16'd5445,-16'd6447,-16'd4041,-16'd6347,-16'd3581,16'd2010,-16'd7472,-16'd1759,16'd3998,-16'd2000,-16'd8771,-16'd4350,16'd6075,16'd4268,16'd6659,16'd5390,-16'd4409,16'd7523,-16'd2667,16'd6941,16'd953,16'd7770,-16'd3810,16'd6129,-16'd2816,-16'd3611,-16'd4540,-16'd4574,16'd3146,-16'd4273};
dout[706]={ -16'd4020,-16'd5902,16'd4956,16'd7233,16'd3312,-16'd1675,-16'd3827,16'd9000,16'd4205,-16'd6008,-16'd2796,-16'd3177,-16'd8107,16'd3156,16'd2154,16'd5050,16'd299,-16'd2290,-16'd750,16'd2977,16'd1268,-16'd1936,-16'd6697,-16'd854,-16'd7942,16'd6088,16'd2731,-16'd2015,-16'd6620,16'd1779,16'd1633,16'd4709,16'd1855,16'd6610,16'd1643,16'd5112};
dout[707]={ -16'd3193,16'd4195,-16'd3251,-16'd7209,16'd4243,16'd3358,-16'd1029,-16'd1140,16'd5919,-16'd6141,16'd2239,16'd541,-16'd4124,16'd1662,16'd3098,-16'd785,-16'd4280,-16'd254,16'd133,-16'd3338,-16'd6554,16'd4630,16'd507,16'd2801,-16'd3261,16'd5149,16'd220,16'd5723,-16'd2011,16'd4097,-16'd2823,-16'd2876,-16'd2462,16'd477,-16'd33,-16'd3188};
dout[708]={ -16'd8485,-16'd6045,16'd3537,-16'd6294,-16'd5347,-16'd266,16'd2830,16'd7809,16'd6498,16'd522,16'd3354,16'd8101,-16'd7645,16'd1061,16'd6504,-16'd1681,-16'd1109,-16'd5192,16'd6314,-16'd53,-16'd4397,-16'd6606,16'd4604,-16'd2096,16'd4895,16'd1926,16'd3543,16'd6669,-16'd3044,16'd3113,16'd2173,16'd4206,16'd7336,-16'd3442,-16'd492,16'd518};
dout[709]={ 16'd5536,16'd2303,-16'd730,16'd939,16'd4712,-16'd4901,-16'd1603,-16'd2324,-16'd1470,16'd4972,-16'd908,-16'd3456,-16'd3493,16'd5788,16'd5357,-16'd3261,16'd5968,16'd3104,-16'd3847,16'd5138,-16'd2769,16'd917,16'd1439,16'd6462,16'd3921,16'd5638,-16'd853,-16'd3697,16'd2146,16'd2979,-16'd2879,16'd3828,-16'd7606,-16'd1151,-16'd1852,16'd3972};
dout[710]={ -16'd7823,16'd8807,16'd3101,-16'd5395,-16'd5676,16'd2082,-16'd19,16'd8656,16'd3607,-16'd3960,-16'd8365,16'd4022,16'd1199,-16'd3488,16'd6682,16'd11813,-16'd6185,-16'd1916,-16'd4648,-16'd9978,16'd6930,-16'd2163,16'd5915,16'd247,-16'd786,16'd3858,-16'd3768,-16'd3111,-16'd9845,-16'd2500,16'd5689,16'd8182,-16'd1089,16'd2745,-16'd7823,16'd7277};
dout[711]={ 16'd2014,16'd3055,-16'd3048,-16'd1771,16'd2747,-16'd1228,16'd2034,16'd5534,16'd554,16'd682,-16'd2586,-16'd4055,-16'd9,16'd4329,-16'd3951,16'd1759,-16'd3655,16'd2909,16'd4985,-16'd6323,16'd2890,16'd4410,16'd1525,16'd1927,-16'd6198,-16'd7747,-16'd6166,16'd4697,16'd237,-16'd3424,-16'd6022,16'd620,-16'd5019,16'd2183,16'd8031,16'd691};
dout[712]={ -16'd2446,16'd4213,16'd2599,-16'd2352,16'd5739,-16'd6138,-16'd963,-16'd3645,16'd6782,-16'd4000,-16'd3306,-16'd7547,-16'd5634,-16'd7730,16'd3114,-16'd3324,-16'd5276,16'd3235,16'd4932,-16'd1794,16'd4466,-16'd2830,-16'd3389,-16'd3021,-16'd6772,16'd1874,16'd0,-16'd5970,-16'd4394,-16'd9151,16'd2953,-16'd8810,-16'd473,-16'd6537,16'd6063,-16'd3189};
dout[713]={ -16'd2016,16'd1066,-16'd2679,16'd864,16'd5575,-16'd2405,16'd2523,-16'd1956,16'd516,16'd829,16'd11673,16'd5783,16'd8443,-16'd4784,16'd2034,16'd783,16'd4347,16'd3770,16'd5673,-16'd6120,16'd308,16'd839,-16'd8375,-16'd3642,16'd3880,-16'd6511,-16'd4082,-16'd12598,-16'd3021,-16'd3222,16'd6796,-16'd7217,-16'd7570,-16'd8119,16'd841,16'd8942};
dout[714]={ 16'd2582,16'd2178,-16'd3937,16'd7222,-16'd1073,16'd7044,-16'd5337,-16'd7230,-16'd6060,-16'd7038,-16'd2218,-16'd7984,-16'd6139,16'd1449,16'd5905,16'd8256,-16'd2297,-16'd7258,16'd3405,16'd1529,-16'd4724,16'd713,16'd272,-16'd4644,-16'd1230,16'd5181,16'd7514,16'd1486,16'd6621,-16'd819,-16'd3495,16'd5468,-16'd7209,-16'd5445,16'd4890,16'd4821};
dout[715]={ -16'd6325,16'd5302,16'd8103,16'd1084,16'd4086,-16'd879,16'd6007,16'd3429,16'd723,16'd3164,16'd5976,-16'd2187,16'd5682,16'd2021,16'd3262,16'd3788,16'd3633,-16'd6734,16'd3449,-16'd7285,16'd7160,16'd4405,-16'd5928,-16'd4982,16'd2056,-16'd5236,-16'd8095,16'd5405,16'd3101,-16'd4407,-16'd3028,16'd8974,-16'd6938,-16'd7451,-16'd1014,16'd2353};
dout[716]={ 16'd1007,-16'd1217,16'd6362,-16'd243,16'd2737,-16'd6512,-16'd1542,-16'd4183,-16'd1735,16'd3813,-16'd776,16'd5321,-16'd2057,-16'd5267,-16'd1916,16'd468,16'd1772,16'd3195,16'd6224,-16'd1871,16'd1501,16'd1892,16'd5233,-16'd764,-16'd6095,16'd1141,16'd662,16'd2804,-16'd420,-16'd1548,16'd2919,16'd370,-16'd3246,-16'd1230,16'd6943,16'd1247};
dout[717]={ -16'd5107,16'd5650,16'd6853,-16'd7691,16'd3808,16'd3526,-16'd3367,16'd2747,-16'd4038,16'd2024,-16'd3872,16'd546,16'd2359,-16'd3324,-16'd2759,-16'd762,16'd1543,-16'd2824,-16'd236,16'd4020,-16'd355,-16'd6174,16'd2942,16'd1630,-16'd6205,16'd2630,-16'd7815,-16'd3877,16'd2217,-16'd7987,16'd4435,16'd5884,-16'd3097,16'd617,16'd2410,-16'd1567};
dout[718]={ -16'd3402,-16'd5131,-16'd1671,-16'd8725,-16'd5549,-16'd2539,16'd5361,-16'd5114,16'd609,16'd5357,16'd6539,-16'd2687,16'd5037,16'd6730,16'd2915,-16'd3127,-16'd3665,16'd5460,-16'd5670,-16'd2326,16'd6236,16'd4960,-16'd7598,16'd4279,16'd6846,-16'd6844,-16'd5649,16'd857,16'd409,-16'd6712,16'd2794,-16'd1473,-16'd1153,-16'd7117,-16'd2561,-16'd2573};
dout[719]={ 16'd3170,16'd5002,-16'd7754,16'd2159,-16'd78,16'd1099,-16'd2849,-16'd4276,16'd4479,16'd4079,-16'd2887,16'd5746,-16'd3763,-16'd1141,16'd1709,16'd6254,16'd6086,16'd2039,16'd4704,-16'd1662,-16'd4003,-16'd6708,-16'd1537,-16'd2923,-16'd3332,16'd6799,16'd2220,-16'd2522,16'd5116,-16'd6187,16'd2846,-16'd5935,-16'd516,16'd4800,16'd5486,-16'd3048};
dout[720]={ -16'd1293,16'd2277,-16'd3759,-16'd3599,-16'd11104,-16'd350,16'd269,-16'd476,-16'd3169,-16'd2172,16'd5177,-16'd5469,16'd2624,16'd143,-16'd2061,16'd6769,16'd2218,16'd2574,-16'd2685,-16'd1461,-16'd8155,-16'd9029,-16'd1425,16'd4753,16'd2872,-16'd9542,16'd8304,16'd7185,-16'd157,16'd5191,16'd3889,16'd3398,-16'd9755,16'd1532,16'd4130,16'd2607};
dout[721]={ 16'd7198,-16'd2540,-16'd1147,16'd4998,16'd4824,-16'd6873,16'd1205,16'd2662,16'd3123,16'd5905,-16'd4127,-16'd4778,16'd3297,16'd3716,-16'd1119,16'd3724,-16'd4865,-16'd5470,16'd2348,-16'd8927,-16'd997,16'd4454,16'd5449,16'd1472,-16'd8846,-16'd1839,-16'd1871,16'd2024,-16'd3102,-16'd5692,-16'd818,-16'd2529,-16'd3203,16'd1136,-16'd6508,16'd6987};
dout[722]={ -16'd886,16'd7881,16'd1018,-16'd269,-16'd3372,16'd6239,-16'd7615,16'd2384,16'd4251,16'd7352,16'd3491,16'd2846,-16'd3886,-16'd11883,-16'd1893,16'd821,16'd1973,-16'd1774,16'd1995,-16'd6307,-16'd5072,16'd3458,-16'd1171,-16'd950,16'd5374,16'd1587,-16'd8985,-16'd6988,16'd2386,-16'd430,-16'd45,16'd890,16'd2933,-16'd912,-16'd4374,16'd188};
dout[723]={ -16'd6294,-16'd2460,16'd3332,-16'd960,16'd572,-16'd1861,-16'd6961,16'd8146,-16'd4221,-16'd6634,16'd8056,-16'd5119,16'd2532,-16'd9137,16'd4776,16'd1184,16'd3086,16'd169,16'd7874,-16'd1188,-16'd7305,16'd3745,-16'd3924,16'd4474,-16'd8038,16'd5415,16'd879,-16'd4136,16'd404,16'd2911,16'd4071,-16'd5464,-16'd7249,-16'd7826,16'd5276,-16'd4930};
dout[724]={ -16'd8805,-16'd5846,16'd4944,16'd2631,16'd3894,16'd807,16'd3579,-16'd5129,-16'd6281,-16'd3046,16'd4956,-16'd5659,16'd7678,16'd822,16'd6111,16'd8490,-16'd4435,-16'd707,-16'd2659,-16'd4229,-16'd11151,16'd5893,16'd1000,16'd2120,-16'd5862,-16'd5398,16'd6115,-16'd9133,-16'd4932,16'd5554,16'd2529,-16'd1779,16'd1713,-16'd6612,16'd3857,16'd4055};
dout[725]={ 16'd2745,16'd2234,16'd5850,16'd3811,-16'd3331,16'd1589,16'd2122,16'd7560,-16'd3380,-16'd1153,-16'd1149,16'd4942,16'd7133,-16'd3506,16'd2612,16'd3102,16'd7167,16'd4619,-16'd3794,-16'd1109,-16'd127,16'd6001,-16'd7346,-16'd1971,16'd1516,-16'd2923,16'd6924,-16'd5685,-16'd447,16'd1035,16'd669,-16'd3331,-16'd7858,16'd262,16'd30,16'd5254};
dout[726]={ 16'd5201,-16'd2991,-16'd4903,-16'd2364,16'd3415,-16'd7299,-16'd1462,-16'd538,-16'd1572,-16'd8489,16'd5172,16'd347,16'd880,16'd1258,-16'd3881,-16'd1435,-16'd5459,16'd2352,16'd6198,16'd4423,-16'd6744,16'd7547,-16'd5424,-16'd4298,16'd2105,16'd3753,16'd1210,16'd2495,16'd2221,-16'd7623,-16'd787,16'd2064,16'd4523,16'd365,16'd1652,-16'd4829};
dout[727]={ 16'd1770,16'd2475,16'd1395,16'd1325,16'd5158,-16'd937,16'd1873,-16'd5822,-16'd3911,16'd2447,16'd5223,-16'd1142,16'd3310,16'd1870,-16'd109,16'd5496,16'd1008,-16'd1224,-16'd5451,16'd4185,16'd5949,-16'd1120,16'd4589,-16'd3612,16'd3911,-16'd2076,-16'd2354,16'd4455,-16'd7295,-16'd2424,16'd5604,-16'd3148,16'd2240,-16'd7148,-16'd3945,16'd988};
dout[728]={ 16'd2825,16'd6135,-16'd820,16'd1984,-16'd5000,-16'd4361,16'd5302,-16'd4641,-16'd2328,-16'd7522,16'd6571,16'd7155,16'd3792,16'd3813,-16'd3467,16'd6765,16'd1329,16'd2531,16'd4734,-16'd2072,-16'd3136,-16'd5554,-16'd6694,-16'd6099,-16'd860,16'd6525,16'd3308,16'd4375,-16'd3395,-16'd7363,-16'd3048,-16'd706,-16'd1970,-16'd169,16'd7438,16'd6429};
dout[729]={ 16'd3096,-16'd452,-16'd296,16'd3809,16'd3692,16'd1984,-16'd768,-16'd2989,16'd1260,-16'd2093,16'd4559,16'd6558,16'd669,16'd4890,-16'd4857,-16'd1892,-16'd5352,-16'd6027,-16'd6039,16'd3256,-16'd4411,-16'd2961,16'd1998,-16'd3734,-16'd5331,-16'd5361,-16'd5013,-16'd4990,-16'd5329,16'd273,16'd5831,16'd4884,-16'd1602,-16'd3839,16'd6611,16'd1705};
dout[730]={ 16'd7468,16'd3253,-16'd2665,-16'd3135,-16'd13197,16'd5014,16'd2189,-16'd1220,16'd5085,-16'd8202,-16'd3023,16'd2268,-16'd1109,-16'd4734,-16'd6457,16'd8768,16'd5527,16'd5430,-16'd121,16'd266,-16'd12773,-16'd3535,16'd6132,16'd5607,-16'd8186,-16'd9632,-16'd890,16'd7317,-16'd9881,16'd4964,16'd2232,-16'd5150,-16'd1748,16'd282,16'd2346,-16'd3176};
dout[731]={ -16'd3869,-16'd1426,-16'd1249,-16'd4688,-16'd6771,-16'd2940,-16'd7731,-16'd5326,-16'd1296,16'd2438,16'd6858,-16'd6477,16'd439,-16'd11098,-16'd2315,16'd68,16'd4740,-16'd7905,16'd1547,-16'd7903,-16'd5628,-16'd4657,-16'd8144,16'd1967,-16'd4590,-16'd6326,-16'd8032,-16'd7714,16'd7464,-16'd1905,-16'd714,-16'd4999,-16'd4029,16'd427,16'd6308,16'd5039};
dout[732]={ 16'd1065,-16'd8277,16'd792,-16'd1404,-16'd2450,16'd3401,-16'd662,16'd5794,16'd2720,16'd7056,-16'd2568,-16'd4836,-16'd9218,-16'd6583,-16'd1701,16'd4497,16'd8940,-16'd2711,-16'd1679,-16'd3984,-16'd2955,-16'd6390,-16'd4912,16'd1693,16'd2766,16'd2026,-16'd6811,-16'd9858,16'd6272,-16'd2489,16'd4881,-16'd3626,16'd2628,-16'd1625,-16'd1490,16'd3325};
dout[733]={ -16'd4981,16'd5773,-16'd834,16'd3134,16'd5790,16'd4442,-16'd6800,16'd3430,16'd3248,-16'd6473,16'd5105,-16'd11758,-16'd7102,16'd546,-16'd2439,16'd3853,16'd2756,-16'd1983,16'd2342,-16'd7482,-16'd8346,16'd3378,-16'd628,-16'd6888,-16'd511,16'd2911,16'd4012,-16'd10908,16'd5108,-16'd849,-16'd3114,-16'd7439,-16'd2146,-16'd7818,16'd8052,-16'd6835};
dout[734]={ 16'd3143,16'd6247,16'd3346,16'd1550,16'd1587,-16'd6336,16'd723,-16'd586,-16'd5757,-16'd5703,16'd4465,-16'd857,16'd8068,-16'd9197,-16'd6542,16'd1008,-16'd4438,-16'd3747,16'd1955,-16'd9926,-16'd11416,16'd4904,-16'd104,16'd5040,-16'd2845,16'd3017,16'd4054,-16'd8433,16'd3404,-16'd4602,16'd5694,16'd232,-16'd2384,16'd4979,16'd6314,-16'd610};
dout[735]={ 16'd995,16'd2734,-16'd2382,-16'd3637,16'd8142,16'd2738,16'd5459,-16'd239,-16'd1425,16'd4743,16'd2145,-16'd2756,16'd7633,-16'd8929,-16'd2564,16'd5924,-16'd317,16'd3093,-16'd2065,16'd5986,-16'd3318,-16'd1347,-16'd5379,16'd1759,16'd3858,16'd7939,-16'd2546,-16'd2777,-16'd5391,-16'd5397,16'd6184,-16'd1017,-16'd4743,16'd2745,-16'd2633,-16'd2182};
dout[736]={ -16'd1855,-16'd7777,-16'd3700,16'd2179,-16'd2833,16'd274,-16'd5605,-16'd4576,16'd5921,16'd3471,-16'd6383,-16'd2516,16'd748,16'd6016,-16'd965,16'd6814,16'd6516,16'd2375,-16'd3172,16'd4343,16'd1434,-16'd4219,-16'd1259,16'd4040,16'd2966,16'd6074,-16'd2352,16'd4924,16'd5561,-16'd6530,-16'd6232,16'd980,16'd494,-16'd3426,-16'd3887,16'd801};
dout[737]={ 16'd496,16'd2520,16'd6905,16'd168,-16'd3327,-16'd4741,-16'd2183,16'd1465,16'd5968,16'd1224,16'd4350,16'd3811,16'd4736,16'd686,16'd1891,-16'd2370,-16'd1322,-16'd8004,-16'd4276,-16'd5570,16'd3142,16'd5289,-16'd3721,-16'd5811,16'd266,-16'd2177,16'd3528,-16'd4392,-16'd5906,-16'd1837,16'd4709,-16'd6382,16'd2222,-16'd7734,-16'd3112,-16'd5122};
dout[738]={ -16'd5802,-16'd5635,-16'd1462,16'd714,16'd4358,16'd6082,16'd5865,-16'd1598,16'd8059,16'd6311,-16'd3578,-16'd3984,16'd1167,16'd6667,16'd2213,16'd6550,16'd5359,-16'd3036,-16'd9369,16'd3343,-16'd7733,-16'd1571,-16'd7591,16'd3029,-16'd2211,-16'd2635,-16'd64,-16'd1209,16'd4285,-16'd3400,16'd1472,-16'd4748,16'd3967,-16'd7072,16'd3095,16'd6163};
dout[739]={ -16'd1893,16'd2069,-16'd1658,-16'd2592,16'd815,16'd5414,-16'd1556,16'd5031,-16'd2157,16'd225,16'd2087,16'd3399,-16'd6693,-16'd5722,-16'd925,-16'd4052,16'd2381,-16'd3548,-16'd9185,-16'd6366,16'd2214,-16'd2854,16'd35,16'd2323,16'd5252,16'd7388,-16'd4244,-16'd7004,16'd1880,-16'd3538,16'd7251,-16'd3680,16'd4168,-16'd1895,16'd3809,16'd4824};
dout[740]={ 16'd7020,16'd1292,16'd92,-16'd6421,-16'd12233,-16'd1448,-16'd9799,-16'd5278,-16'd5494,-16'd7127,-16'd465,16'd2745,-16'd2702,-16'd7326,-16'd1113,16'd1609,16'd10964,-16'd1050,16'd207,16'd11957,-16'd13979,-16'd11073,-16'd6287,16'd453,16'd5599,-16'd10356,16'd381,-16'd1456,-16'd3239,-16'd3340,16'd4718,-16'd391,16'd3990,-16'd8997,-16'd2476,16'd1903};
dout[741]={ 16'd1607,-16'd4579,-16'd1718,-16'd1370,16'd2385,16'd4383,16'd4029,16'd190,16'd2607,-16'd1247,16'd11350,-16'd6044,-16'd3517,16'd5043,-16'd12522,16'd3800,16'd7750,16'd4234,-16'd7330,16'd2521,-16'd5851,16'd3662,-16'd8315,16'd6964,16'd3536,-16'd7284,16'd1628,16'd2441,-16'd1442,-16'd2670,-16'd1657,-16'd9028,-16'd7655,-16'd8495,-16'd8893,-16'd5202};
dout[742]={ -16'd7693,-16'd167,16'd592,16'd8859,16'd3859,-16'd7822,16'd316,16'd7161,16'd6184,-16'd7393,16'd9200,-16'd9747,-16'd9484,-16'd8334,-16'd7411,16'd2625,16'd1419,16'd237,-16'd6276,-16'd6794,-16'd5369,16'd4331,-16'd2860,-16'd6974,16'd5544,-16'd10565,-16'd1438,16'd2321,-16'd558,-16'd5779,-16'd4896,-16'd4332,-16'd5228,-16'd6363,16'd3032,-16'd4628};
dout[743]={ -16'd1824,-16'd5471,16'd2423,16'd3016,-16'd2342,-16'd5396,-16'd8859,16'd7427,16'd2588,16'd3399,16'd8501,-16'd8726,16'd1772,-16'd7455,-16'd1735,16'd3530,-16'd3197,-16'd1454,16'd789,-16'd1781,-16'd624,16'd372,-16'd280,16'd3868,-16'd6524,16'd6731,16'd7218,-16'd7778,16'd3840,16'd8140,16'd3256,-16'd4932,-16'd5853,-16'd3415,-16'd1173,16'd2417};
dout[744]={ 16'd3356,-16'd80,16'd2115,16'd6375,16'd3912,-16'd4638,-16'd5597,16'd3790,-16'd7005,-16'd8553,-16'd1197,16'd4910,-16'd3791,-16'd9375,-16'd7080,-16'd1770,-16'd6302,16'd3877,16'd7379,16'd2927,-16'd2071,-16'd90,-16'd6193,16'd1920,16'd6792,16'd2026,16'd288,-16'd3709,16'd1667,16'd1197,-16'd653,-16'd2847,-16'd785,16'd114,16'd2421,-16'd2106};
dout[745]={ -16'd6404,-16'd5909,16'd2516,-16'd6454,-16'd747,-16'd6425,-16'd4507,-16'd4170,-16'd1125,-16'd2310,-16'd5695,16'd642,16'd3766,16'd3386,16'd4233,-16'd4551,-16'd5681,16'd6237,-16'd5462,-16'd5715,-16'd1960,16'd4054,-16'd374,16'd2713,-16'd1390,-16'd2124,-16'd1318,-16'd5370,-16'd3131,16'd895,-16'd475,-16'd6897,-16'd4130,-16'd2228,-16'd2819,16'd9346};
dout[746]={ 16'd6052,-16'd6939,16'd1557,16'd2546,-16'd3476,-16'd5607,-16'd6943,16'd2795,-16'd5833,16'd5047,16'd1523,16'd2166,16'd6996,16'd4801,-16'd2035,16'd6511,16'd5594,-16'd7748,-16'd681,-16'd4513,-16'd7422,16'd4835,16'd5312,16'd6435,16'd90,-16'd3408,16'd3508,16'd3577,16'd6423,16'd4057,16'd7828,-16'd8828,16'd4539,-16'd3833,-16'd2836,16'd2416};
dout[747]={ 16'd4495,-16'd1750,-16'd318,16'd1336,16'd549,-16'd6111,16'd3273,-16'd4767,16'd3826,16'd10,16'd701,16'd4340,16'd4141,16'd3985,-16'd3130,-16'd3303,16'd7320,-16'd8630,16'd2274,16'd4668,16'd1663,16'd3892,16'd1393,-16'd30,-16'd8603,16'd7960,-16'd4265,16'd4381,16'd8494,16'd5879,-16'd2756,16'd2442,-16'd407,-16'd3610,-16'd5601,16'd6351};
dout[748]={ -16'd986,16'd6249,16'd3876,-16'd6851,-16'd598,16'd5010,16'd207,-16'd2596,16'd4119,-16'd3214,16'd4150,16'd1123,-16'd457,16'd4829,-16'd2115,16'd4142,16'd5254,16'd2272,-16'd9658,-16'd4571,16'd3625,-16'd1351,16'd5718,16'd161,-16'd4371,16'd753,-16'd4582,16'd6531,-16'd3951,-16'd3938,16'd972,16'd4582,16'd3770,-16'd2568,-16'd5936,16'd2725};
dout[749]={ 16'd5365,16'd2412,-16'd6116,-16'd1558,-16'd3547,16'd2569,-16'd3818,-16'd343,16'd6408,-16'd650,-16'd2680,16'd5767,-16'd684,16'd8051,-16'd1568,16'd4452,16'd2512,-16'd4510,-16'd7532,16'd2616,-16'd4995,-16'd5861,16'd5197,16'd2608,16'd4405,16'd831,16'd573,-16'd3692,16'd4870,-16'd6399,16'd1040,-16'd954,16'd4347,-16'd2538,16'd2979,-16'd6900};
dout[750]={ -16'd3340,-16'd5154,-16'd5644,-16'd1247,-16'd13757,16'd4221,-16'd1674,-16'd5901,-16'd3350,16'd4658,16'd724,16'd1359,-16'd4049,-16'd4265,-16'd732,-16'd358,16'd3286,-16'd1833,-16'd9134,16'd3590,16'd275,-16'd422,16'd5419,-16'd1366,-16'd5375,-16'd8216,16'd6873,-16'd5721,16'd1188,-16'd4157,16'd6395,16'd1946,-16'd3363,16'd3872,-16'd5153,-16'd3466};
dout[751]={ -16'd6037,-16'd5936,16'd4032,-16'd2922,16'd5349,-16'd4974,-16'd5587,16'd2413,16'd2954,-16'd7013,16'd12118,16'd217,-16'd7782,-16'd4582,-16'd2691,16'd1072,-16'd7238,16'd34,16'd3468,16'd6515,-16'd4408,-16'd4801,16'd2195,16'd6167,16'd578,-16'd674,-16'd122,16'd4115,16'd7319,-16'd7063,-16'd3117,-16'd2581,16'd2052,-16'd5099,-16'd13206,-16'd5044};
dout[752]={ -16'd5526,-16'd2919,16'd2217,16'd9228,-16'd3618,-16'd4815,16'd473,-16'd4176,-16'd5368,16'd1538,16'd9720,-16'd4655,-16'd7653,-16'd2398,-16'd3797,-16'd318,16'd4676,16'd6856,16'd5780,16'd4947,-16'd3064,16'd1859,-16'd3,16'd4630,-16'd5085,-16'd2371,-16'd2320,16'd1286,-16'd1021,16'd5570,-16'd4988,-16'd9266,-16'd740,16'd3012,-16'd12877,16'd974};
dout[753]={ -16'd819,16'd7858,16'd3157,-16'd401,-16'd2807,-16'd4100,-16'd6673,16'd8320,16'd3302,16'd3828,-16'd7842,-16'd5276,-16'd10785,16'd2047,-16'd4613,-16'd896,-16'd1037,16'd588,16'd7943,-16'd1819,16'd4186,16'd2156,16'd5142,16'd9113,16'd3858,-16'd6957,16'd476,-16'd8316,-16'd2330,16'd5288,-16'd7283,16'd2400,-16'd8787,16'd836,16'd73,16'd1695};
dout[754]={ -16'd7036,16'd6520,-16'd2662,-16'd9159,-16'd2194,-16'd3937,16'd1236,-16'd4899,16'd2487,16'd527,-16'd4122,16'd140,-16'd7558,-16'd9865,-16'd428,16'd2668,-16'd3383,16'd5892,16'd4191,16'd639,16'd7372,16'd1569,-16'd4042,-16'd2742,-16'd1851,16'd1984,16'd6036,16'd1840,16'd1176,-16'd1367,16'd1107,-16'd9627,-16'd16,-16'd2400,-16'd2575,-16'd1515};
dout[755]={ -16'd8632,16'd2661,-16'd2000,-16'd6686,-16'd915,-16'd5269,16'd1416,16'd1513,16'd1235,16'd108,16'd1619,16'd4776,16'd4695,-16'd1720,16'd1704,-16'd4106,-16'd4925,-16'd3634,-16'd5989,16'd2391,-16'd1751,-16'd588,16'd1987,-16'd3418,-16'd5770,16'd2477,16'd113,16'd1891,-16'd3389,16'd4485,-16'd5111,-16'd3074,16'd1307,16'd5057,-16'd903,16'd4757};
dout[756]={ -16'd2135,-16'd6209,16'd4204,16'd2387,-16'd3106,16'd2085,-16'd3671,16'd540,-16'd4425,16'd6774,16'd7730,-16'd3460,-16'd8202,-16'd7952,16'd3202,16'd5734,-16'd7715,16'd1619,-16'd2296,16'd2514,16'd949,16'd2832,-16'd3624,-16'd4136,16'd548,16'd304,16'd5079,-16'd6037,-16'd3059,-16'd3760,-16'd5449,-16'd1678,-16'd1537,16'd3773,-16'd2603,-16'd3086};
dout[757]={ 16'd3680,-16'd5709,-16'd7591,16'd692,-16'd2572,16'd3416,16'd4558,16'd5930,-16'd470,-16'd235,16'd2120,16'd6640,-16'd973,16'd487,16'd5281,-16'd4799,-16'd4421,-16'd2151,16'd2497,16'd2960,16'd7326,-16'd5367,-16'd5667,-16'd7489,-16'd5183,-16'd4587,-16'd1528,-16'd7508,16'd3723,-16'd167,16'd4403,16'd2456,16'd5852,16'd933,-16'd2174,16'd2812};
dout[758]={ 16'd2541,-16'd776,16'd3843,-16'd7102,16'd7331,16'd856,-16'd4379,-16'd2682,-16'd561,-16'd4833,16'd5517,-16'd4401,16'd2249,16'd5163,16'd1716,-16'd4730,-16'd4869,16'd5108,-16'd9231,16'd3786,-16'd2076,16'd3547,16'd3978,-16'd8790,-16'd2115,16'd1213,16'd2930,-16'd3794,-16'd6161,-16'd4388,16'd5501,-16'd4270,-16'd1305,-16'd9195,-16'd4330,-16'd1150};
dout[759]={ -16'd5743,-16'd1862,-16'd3654,16'd4950,-16'd5694,-16'd5547,-16'd101,16'd326,16'd474,-16'd3384,-16'd3528,16'd4572,16'd2142,16'd4935,16'd2206,16'd4588,16'd1101,16'd5619,-16'd2524,-16'd2613,-16'd5997,16'd3017,16'd3556,-16'd2149,16'd9,-16'd2572,16'd4691,16'd4240,-16'd2869,16'd3571,16'd6659,-16'd8281,-16'd4713,-16'd8103,-16'd3627,-16'd5823};
dout[760]={ 16'd6097,-16'd8523,-16'd592,-16'd860,-16'd4681,-16'd2111,-16'd1212,16'd1337,-16'd3544,-16'd1577,16'd9384,16'd7884,-16'd5652,16'd7360,-16'd4211,16'd2481,16'd5154,-16'd6877,16'd3375,16'd4915,16'd5849,16'd7584,-16'd5517,-16'd6976,-16'd8651,16'd1273,16'd4898,-16'd2557,-16'd7629,-16'd4042,16'd2732,-16'd3752,-16'd2653,16'd6727,-16'd8628,16'd5237};
dout[761]={ 16'd2926,16'd6158,-16'd3037,16'd1709,16'd2030,16'd2103,-16'd5194,-16'd4472,16'd1989,16'd5508,16'd4087,16'd7600,16'd2203,16'd2449,-16'd4796,16'd7224,-16'd7004,-16'd5054,16'd3453,16'd1519,16'd4355,-16'd4070,-16'd3156,-16'd18,16'd799,16'd5661,16'd4298,-16'd5671,-16'd6509,-16'd8148,-16'd7587,-16'd992,-16'd4080,-16'd3769,-16'd10467,-16'd796};
dout[762]={ -16'd7304,-16'd6080,16'd5765,16'd5283,-16'd6338,16'd1579,16'd6046,-16'd7334,16'd2978,16'd4628,16'd4913,-16'd352,-16'd4338,16'd7755,16'd1289,16'd5416,-16'd5159,16'd4690,-16'd493,-16'd3553,16'd7597,16'd7504,-16'd4491,16'd1832,-16'd3026,-16'd7049,16'd6657,16'd3001,-16'd4149,-16'd3419,-16'd7694,-16'd3435,-16'd6095,-16'd5971,-16'd6163,-16'd4747};
dout[763]={ 16'd3770,-16'd1565,-16'd2311,16'd1537,16'd825,-16'd3062,16'd1333,-16'd6019,16'd4649,-16'd577,16'd1957,-16'd629,-16'd10673,16'd2169,-16'd6909,16'd1833,-16'd4199,-16'd3339,-16'd2159,-16'd1513,16'd2253,16'd2419,-16'd2383,16'd7953,16'd1160,16'd1583,16'd8101,16'd4126,16'd4008,-16'd4920,-16'd2178,-16'd5396,-16'd6824,-16'd2654,-16'd1331,-16'd6079};
dout[764]={ -16'd8670,-16'd5033,16'd1526,16'd1897,16'd8513,16'd186,-16'd5222,-16'd135,16'd3494,-16'd5423,16'd47,16'd1460,-16'd5351,-16'd7707,-16'd5068,16'd1494,-16'd4959,16'd5171,16'd1151,16'd3418,16'd6285,16'd4423,-16'd5663,16'd7147,-16'd3454,16'd2000,-16'd1861,-16'd6979,16'd3459,16'd6266,-16'd5580,16'd538,-16'd3646,-16'd3190,16'd3378,16'd7109};
dout[765]={ 16'd2489,16'd5266,16'd1755,-16'd4674,16'd7323,-16'd4211,16'd2738,16'd6704,-16'd207,-16'd4123,16'd5091,16'd4351,-16'd4190,-16'd5424,-16'd1069,-16'd8586,-16'd7406,16'd3541,16'd988,16'd3382,-16'd2710,16'd3079,16'd4478,-16'd4965,-16'd7590,-16'd2505,16'd4678,-16'd8667,-16'd4859,-16'd5194,-16'd138,-16'd6697,-16'd1703,-16'd1310,16'd6548,-16'd2623};
dout[766]={ -16'd5033,-16'd7784,16'd2787,16'd2994,-16'd5648,16'd4347,-16'd2261,16'd1024,-16'd1600,16'd1549,-16'd1705,16'd6035,-16'd4601,-16'd7723,16'd1327,-16'd3020,-16'd7229,-16'd1834,-16'd3191,16'd1440,-16'd5202,16'd4243,16'd3989,-16'd6457,16'd5642,-16'd3631,-16'd4352,-16'd1519,16'd699,16'd5525,16'd2245,-16'd5015,-16'd1877,16'd1821,-16'd6829,16'd666};
dout[767]={ 16'd468,16'd5295,-16'd7156,16'd6253,-16'd987,-16'd2443,-16'd6439,-16'd2753,16'd3269,-16'd704,-16'd2294,16'd3031,-16'd799,16'd7175,-16'd2779,16'd4297,-16'd8773,16'd2996,-16'd5898,16'd675,-16'd6056,16'd83,16'd6446,-16'd7571,-16'd5287,-16'd3205,-16'd5238,-16'd7266,-16'd1660,16'd824,16'd2392,16'd7001,16'd153,16'd3472,16'd5332,16'd2056};
dout[768]={ -16'd3750,-16'd4310,16'd2524,16'd1057,-16'd108,16'd5032,-16'd7455,-16'd6107,16'd5424,16'd1823,-16'd4924,16'd4260,-16'd4847,-16'd1627,-16'd4867,-16'd2931,-16'd6421,16'd2704,-16'd4746,16'd3704,16'd953,-16'd5801,-16'd5479,-16'd7737,16'd7766,16'd1603,16'd152,-16'd8294,16'd3358,16'd2311,-16'd6688,16'd2905,16'd5396,16'd1355,16'd2229,-16'd2569};
dout[769]={ -16'd906,-16'd3997,16'd3771,16'd5204,16'd1878,16'd1227,-16'd7051,-16'd614,16'd1853,-16'd2169,-16'd4774,16'd6260,-16'd6010,16'd5792,16'd9782,-16'd5568,-16'd4713,-16'd1735,-16'd7209,-16'd5267,16'd58,16'd5492,16'd5223,-16'd8809,16'd2497,16'd787,16'd1660,-16'd5092,16'd6532,16'd1356,-16'd7213,16'd4698,16'd4779,16'd3529,-16'd8355,-16'd10514};
dout[770]={ 16'd2725,-16'd8581,-16'd2974,16'd3548,-16'd8236,-16'd7877,-16'd9496,-16'd1427,16'd3025,-16'd4799,16'd10463,-16'd4032,16'd3089,-16'd3186,16'd2701,-16'd6685,-16'd5207,-16'd7106,16'd7481,16'd3200,-16'd2550,16'd7915,16'd4540,16'd3190,-16'd9147,16'd3364,16'd7506,-16'd8120,-16'd6983,-16'd348,16'd628,-16'd7443,-16'd6846,-16'd3562,-16'd12017,16'd3640};
dout[771]={ 16'd8011,16'd4907,-16'd1742,-16'd2955,-16'd2869,-16'd4989,-16'd6716,16'd702,-16'd7673,-16'd3607,-16'd791,16'd2876,-16'd1696,-16'd1766,-16'd8211,16'd3494,-16'd5673,-16'd2343,-16'd3003,16'd4705,-16'd6510,16'd441,-16'd7041,-16'd4122,16'd4215,16'd7986,16'd3050,16'd5768,-16'd8445,-16'd3998,-16'd9606,16'd4934,-16'd7191,-16'd5649,-16'd9281,-16'd5182};
dout[772]={ -16'd8549,-16'd4043,16'd938,16'd9098,-16'd2478,-16'd4593,-16'd1182,-16'd4072,16'd5418,16'd1845,-16'd866,16'd7060,-16'd6577,-16'd218,-16'd7115,16'd4977,-16'd10932,16'd1022,-16'd7170,-16'd5054,16'd913,16'd6387,16'd1113,-16'd7205,-16'd3669,-16'd2411,16'd3043,16'd1506,-16'd6183,-16'd8140,-16'd9740,-16'd2926,16'd3515,-16'd951,-16'd12318,-16'd5935};
dout[773]={ 16'd2730,16'd2087,-16'd3705,-16'd6532,-16'd2366,-16'd815,-16'd6262,-16'd6827,-16'd4938,-16'd3660,-16'd4229,-16'd2206,-16'd9582,-16'd2132,16'd5113,-16'd1605,-16'd514,-16'd1790,16'd3719,16'd10609,16'd4785,-16'd1823,-16'd7206,16'd8061,16'd3642,-16'd14174,16'd4662,-16'd4021,-16'd6179,16'd1418,-16'd807,-16'd1268,-16'd7414,16'd5679,16'd2871,16'd4203};
dout[774]={ -16'd6829,-16'd4475,-16'd3547,16'd2420,-16'd563,-16'd2422,-16'd1588,-16'd3352,16'd1678,-16'd181,16'd3712,-16'd2914,-16'd9137,16'd1197,-16'd2231,-16'd6132,-16'd10586,16'd81,-16'd4471,16'd9921,-16'd4393,-16'd1483,-16'd7782,16'd6587,16'd5286,-16'd5177,16'd963,-16'd1841,-16'd5423,16'd1774,16'd1160,16'd473,-16'd9031,16'd1910,-16'd9312,-16'd4553};
dout[775]={ -16'd6905,16'd5507,16'd667,-16'd7291,-16'd4304,-16'd5126,-16'd36,16'd4767,16'd9678,16'd4825,-16'd6089,16'd2,-16'd4523,-16'd3,-16'd8631,-16'd5543,-16'd3569,16'd912,-16'd3808,16'd2980,16'd7717,-16'd3040,-16'd7077,16'd224,16'd277,16'd2812,16'd100,16'd1025,-16'd6645,16'd1108,-16'd8878,-16'd1479,-16'd7384,16'd3681,-16'd366,-16'd1263};
dout[776]={ -16'd8749,16'd4376,-16'd3456,16'd2831,16'd1736,16'd4530,16'd4897,16'd5049,-16'd2354,-16'd2316,16'd741,-16'd1383,-16'd4555,-16'd6335,16'd1162,16'd3459,16'd4877,16'd5059,-16'd2240,16'd436,16'd5254,16'd878,16'd5174,-16'd5616,-16'd1659,16'd6312,16'd6067,16'd52,16'd5195,16'd6907,16'd4942,16'd4160,-16'd2733,16'd3407,16'd1954,-16'd4588};
dout[777]={ 16'd899,-16'd6391,-16'd6818,-16'd5490,-16'd3062,-16'd6350,16'd2760,16'd4447,-16'd3948,-16'd5771,-16'd1712,16'd2896,-16'd5757,16'd5445,-16'd3815,16'd3256,16'd1143,-16'd2140,16'd2757,-16'd212,-16'd5750,16'd1898,-16'd1387,-16'd6087,16'd4279,-16'd5214,-16'd6727,16'd3267,-16'd1620,16'd6853,-16'd7721,-16'd5420,-16'd4881,16'd2444,-16'd2275,-16'd2027};
dout[778]={ 16'd3367,-16'd249,-16'd390,-16'd4568,-16'd1404,-16'd5358,16'd6002,-16'd1435,-16'd1408,-16'd4971,-16'd1324,-16'd675,16'd5318,16'd5674,-16'd6473,16'd2212,16'd3949,-16'd2744,16'd863,-16'd6062,16'd3985,-16'd5180,16'd4311,-16'd28,16'd2527,16'd2805,-16'd3199,-16'd7729,16'd810,16'd7619,-16'd4748,-16'd5705,16'd4679,-16'd4000,-16'd3770,-16'd7399};
dout[779]={ -16'd6772,-16'd7275,16'd9084,16'd5441,16'd1614,16'd5035,16'd7577,-16'd3719,16'd1691,-16'd318,-16'd1463,-16'd4155,16'd2351,16'd5160,-16'd4304,16'd4908,-16'd5631,-16'd7889,-16'd2029,-16'd7019,16'd1106,16'd3588,16'd1681,-16'd2309,16'd4355,16'd276,-16'd360,16'd4622,-16'd6392,16'd7563,16'd2627,16'd6429,16'd2074,16'd4954,-16'd5115,-16'd4739};
dout[780]={ -16'd3411,-16'd6641,16'd4302,16'd6960,-16'd1703,-16'd5516,-16'd2939,-16'd5543,-16'd4526,-16'd6893,16'd7106,16'd3711,-16'd6479,16'd7348,16'd1754,-16'd7774,-16'd2537,16'd2925,-16'd6413,-16'd842,-16'd6668,16'd15235,-16'd1408,16'd800,16'd6043,16'd3551,16'd3508,-16'd4538,-16'd1137,16'd1808,16'd2155,16'd3447,-16'd5245,16'd9913,-16'd2210,-16'd6457};
dout[781]={ 16'd1552,-16'd224,-16'd4039,16'd2092,-16'd5172,-16'd6049,16'd4932,-16'd7586,16'd2848,-16'd2069,16'd10303,-16'd2006,-16'd2008,16'd8077,16'd2634,-16'd4260,-16'd7320,-16'd8362,16'd3999,-16'd1595,-16'd6773,16'd10040,16'd5037,16'd1340,-16'd5535,16'd5869,16'd2539,16'd6218,-16'd1039,-16'd13604,-16'd131,16'd2764,-16'd5823,-16'd1331,-16'd263,16'd1153};
dout[782]={ -16'd757,-16'd753,16'd976,16'd2635,16'd4055,-16'd3814,-16'd6244,-16'd5132,16'd2290,-16'd4812,16'd2054,16'd1538,16'd671,16'd3651,16'd2829,16'd7588,-16'd6217,-16'd1930,-16'd6944,-16'd5377,-16'd5076,16'd9667,-16'd6935,-16'd5532,-16'd7379,-16'd7291,16'd4684,-16'd782,-16'd4003,-16'd11845,-16'd1591,-16'd830,16'd5888,-16'd5574,-16'd7494,16'd8016};
dout[783]={ 16'd5937,-16'd2137,16'd1931,16'd7780,16'd4833,-16'd2368,-16'd3847,-16'd8709,16'd5836,-16'd7837,-16'd3225,16'd2562,-16'd4946,-16'd812,16'd4441,16'd318,16'd2304,16'd3762,-16'd3542,16'd1869,16'd5641,16'd4237,-16'd6629,-16'd6654,16'd342,-16'd11634,16'd3235,16'd244,-16'd6517,-16'd9089,-16'd2858,-16'd753,-16'd57,-16'd4118,-16'd1008,16'd2604};
dout[784]={ 16'd3649,16'd509,-16'd5774,16'd512,16'd5245,-16'd5860,-16'd6166,-16'd5029,16'd6346,-16'd2737,-16'd5199,-16'd5188,16'd1171,16'd2455,16'd4095,-16'd2259,-16'd3992,-16'd5806,16'd5134,16'd11105,-16'd1374,-16'd4399,-16'd1144,16'd8024,-16'd5650,-16'd5784,-16'd3009,-16'd8156,16'd271,-16'd4489,-16'd5468,16'd3001,-16'd774,16'd257,-16'd2565,-16'd3078};
dout[785]={ -16'd72,16'd5143,16'd6164,-16'd1901,16'd8302,16'd4647,-16'd3581,16'd5803,16'd999,-16'd560,16'd3748,16'd52,-16'd8002,16'd1263,-16'd7496,16'd3912,16'd5921,16'd5076,-16'd7185,16'd5921,16'd7858,-16'd652,16'd6028,16'd6591,-16'd1568,16'd3777,-16'd7603,-16'd8399,-16'd1461,16'd6422,16'd6953,-16'd8839,-16'd2795,16'd4180,16'd1094,-16'd2206};
dout[786]={ 16'd3466,-16'd4320,-16'd8095,16'd2667,16'd4254,-16'd4413,-16'd6141,-16'd6794,16'd3251,-16'd5979,-16'd1934,-16'd5166,16'd6454,16'd5666,-16'd4716,-16'd4924,16'd5656,-16'd1007,16'd2974,-16'd1417,-16'd6230,16'd6876,-16'd7518,16'd6101,16'd2143,-16'd3239,16'd2838,-16'd5509,-16'd490,-16'd949,16'd227,-16'd6489,-16'd6637,16'd3652,-16'd1541,-16'd4274};
dout[787]={ 16'd3335,-16'd6948,-16'd7644,-16'd2571,-16'd7107,16'd7481,16'd4219,-16'd2952,16'd3898,16'd3132,-16'd6414,-16'd3470,16'd2760,-16'd6331,-16'd1637,-16'd1709,-16'd1110,-16'd5374,-16'd232,16'd3349,16'd6239,16'd3716,16'd7254,-16'd4300,-16'd5355,-16'd3535,16'd277,16'd5155,16'd2930,-16'd3390,-16'd2669,-16'd6129,16'd4228,16'd3134,-16'd6362,16'd4825};
dout[788]={ -16'd6583,-16'd4445,-16'd3499,16'd4732,16'd5799,16'd1764,-16'd6412,16'd319,16'd3897,16'd7072,16'd2022,16'd855,16'd4031,-16'd3086,-16'd732,16'd4050,16'd6741,16'd3169,16'd7624,-16'd1853,-16'd3830,16'd6900,-16'd1136,16'd600,16'd5997,-16'd3474,16'd3804,-16'd8018,16'd3783,-16'd5734,16'd5390,-16'd4824,-16'd3070,16'd3227,16'd4494,-16'd719};
dout[789]={ -16'd1960,16'd3924,16'd6668,-16'd5683,-16'd168,16'd2524,16'd3399,16'd3185,-16'd1624,16'd1560,-16'd592,16'd2477,-16'd5060,-16'd7926,16'd3151,-16'd1373,16'd1914,16'd7135,16'd4440,-16'd6016,16'd6517,-16'd816,16'd82,-16'd4942,-16'd2603,-16'd8966,-16'd2754,16'd4945,16'd6784,-16'd2119,16'd3932,16'd7188,-16'd5174,-16'd887,16'd68,16'd725};
dout[790]={ -16'd5437,16'd2854,-16'd8216,16'd8286,16'd2209,-16'd5925,-16'd2961,-16'd545,-16'd1905,-16'd765,16'd2583,-16'd2036,-16'd775,-16'd4607,-16'd1897,-16'd2099,-16'd96,16'd4092,-16'd5309,16'd6834,-16'd4014,16'd10057,-16'd1109,16'd3643,-16'd332,16'd9589,-16'd5595,16'd2782,16'd481,-16'd1005,-16'd651,-16'd5218,-16'd6416,16'd2021,-16'd3060,16'd1679};
dout[791]={ 16'd70,-16'd2061,-16'd4574,-16'd2189,-16'd392,-16'd3037,16'd872,-16'd2784,-16'd2052,-16'd2987,16'd6799,16'd7845,-16'd5838,16'd1857,16'd5680,16'd8221,16'd2731,16'd4616,16'd2491,-16'd702,16'd3206,16'd7004,16'd1147,16'd1959,16'd1215,16'd4553,16'd7082,16'd3961,-16'd3556,-16'd12742,16'd8263,-16'd7804,-16'd590,16'd52,16'd260,16'd2525};
dout[792]={ 16'd4742,16'd7116,16'd5918,16'd2534,16'd7178,16'd6055,16'd4085,-16'd4432,-16'd4752,16'd487,16'd3018,16'd6990,-16'd8997,16'd5326,-16'd2881,-16'd1600,-16'd3463,-16'd2175,-16'd7375,-16'd7940,16'd642,16'd4560,-16'd3984,-16'd430,-16'd2535,-16'd664,16'd283,-16'd3468,-16'd1725,-16'd7518,16'd313,16'd3476,16'd274,16'd3617,-16'd5897,-16'd4372};
dout[793]={ 16'd4649,-16'd3157,16'd1465,-16'd3151,16'd2498,16'd2271,-16'd1461,16'd1739,-16'd2637,16'd2706,16'd5399,-16'd4231,16'd857,16'd4814,-16'd5702,-16'd177,-16'd1697,-16'd6288,16'd5117,16'd7170,16'd564,-16'd5044,-16'd4104,-16'd8177,-16'd4383,-16'd4303,-16'd1757,-16'd6562,-16'd435,-16'd8693,-16'd2268,-16'd3199,-16'd287,16'd3612,16'd1720,-16'd4374};
dout[794]={ 16'd3414,-16'd4483,16'd4303,16'd1499,-16'd6089,-16'd8798,16'd5508,16'd624,-16'd1169,16'd2401,-16'd2889,16'd814,-16'd5637,-16'd2663,16'd5121,-16'd5807,16'd5858,-16'd6557,16'd3657,16'd1627,16'd2877,-16'd6928,16'd7741,16'd1486,-16'd2968,-16'd773,-16'd4995,16'd2286,16'd377,16'd4376,16'd283,16'd3664,-16'd646,16'd5665,16'd1881,-16'd4271};
dout[795]={ -16'd8130,16'd1803,-16'd5242,16'd7249,16'd1241,16'd233,16'd2887,16'd2673,16'd2347,16'd3705,-16'd133,-16'd8170,16'd7235,-16'd178,16'd1574,16'd2367,16'd3512,-16'd6379,16'd6186,16'd4218,-16'd648,16'd805,16'd2283,16'd7386,-16'd5808,-16'd3869,-16'd6436,-16'd2044,16'd6910,16'd6133,-16'd3595,-16'd5145,-16'd6515,16'd1482,-16'd3722,16'd1916};
dout[796]={ -16'd5032,-16'd9014,-16'd2236,-16'd4740,-16'd6674,16'd3030,16'd5289,16'd5465,16'd4116,-16'd6770,16'd5560,16'd3429,16'd8203,-16'd1757,16'd4706,16'd3389,-16'd3863,-16'd1099,16'd717,-16'd3204,16'd6431,-16'd4736,16'd6243,-16'd1256,-16'd5608,-16'd318,-16'd5683,-16'd7126,-16'd3342,16'd6448,-16'd4497,16'd4412,16'd3653,16'd1450,16'd8646,16'd2984};
dout[797]={ 16'd906,16'd346,16'd438,16'd5195,16'd419,16'd4106,-16'd3187,16'd3741,16'd2547,-16'd3697,16'd72,-16'd6522,-16'd3690,16'd5703,16'd3050,16'd4747,-16'd3574,-16'd6576,-16'd1846,-16'd172,-16'd2881,16'd6125,16'd415,16'd4073,16'd589,16'd1264,16'd4782,-16'd4381,16'd2902,-16'd1057,-16'd6833,16'd4127,16'd4072,-16'd7447,-16'd4655,-16'd4339};
dout[798]={ -16'd8769,-16'd6575,16'd3650,16'd10,16'd2472,16'd6797,-16'd3066,16'd2790,-16'd935,-16'd1703,-16'd2650,-16'd5710,-16'd3345,16'd3782,-16'd4878,16'd2327,-16'd479,16'd2842,-16'd1434,-16'd68,-16'd4353,-16'd1195,16'd5062,16'd1232,16'd345,-16'd4301,-16'd5972,-16'd5028,16'd2498,-16'd5852,-16'd5962,-16'd5735,16'd4451,16'd4598,16'd77,16'd1617};
dout[799]={ -16'd6985,16'd1489,16'd2932,-16'd696,-16'd4516,16'd6991,-16'd3370,-16'd156,16'd5947,16'd3493,-16'd4897,-16'd2220,16'd6800,-16'd6229,-16'd5756,16'd2814,16'd2829,16'd764,16'd2180,-16'd3837,16'd5987,16'd5395,16'd118,16'd70,-16'd7637,16'd2631,16'd6355,-16'd5361,-16'd6322,16'd1369,16'd3682,16'd11,-16'd5433,-16'd6428,16'd3287,16'd3363};
dout[800]={ -16'd4894,-16'd2198,-16'd1775,-16'd1814,-16'd7266,-16'd11083,-16'd6961,16'd6296,-16'd8190,-16'd3844,16'd9281,-16'd6173,-16'd4314,16'd4686,-16'd3537,-16'd6397,16'd6041,-16'd1602,-16'd1034,-16'd7310,16'd2014,16'd11467,-16'd1588,-16'd1523,16'd4345,16'd7962,-16'd826,16'd4470,16'd567,16'd3249,-16'd5158,16'd558,-16'd3729,-16'd4194,-16'd10200,-16'd1682};
dout[801]={ -16'd869,-16'd9016,-16'd3060,-16'd2718,-16'd2725,-16'd820,-16'd3664,16'd5035,-16'd7973,-16'd8037,16'd1210,16'd3802,16'd6124,16'd5312,-16'd5699,16'd3455,-16'd1187,-16'd2964,16'd4475,16'd5341,-16'd306,16'd4819,-16'd2319,-16'd3042,-16'd7545,-16'd6321,-16'd2863,16'd5153,-16'd8189,-16'd1107,16'd3772,-16'd7147,16'd5562,-16'd7021,16'd3822,16'd353};
dout[802]={ 16'd5727,16'd5497,-16'd1063,16'd4270,-16'd5556,-16'd2257,-16'd7183,-16'd7021,-16'd6476,16'd3817,-16'd1004,16'd1523,-16'd7372,-16'd26,-16'd3414,16'd8289,-16'd732,-16'd6724,16'd4197,-16'd2704,16'd3074,-16'd7118,-16'd6657,-16'd8190,-16'd8006,16'd2910,-16'd381,-16'd79,16'd452,-16'd8046,16'd3412,16'd2517,-16'd7311,16'd1093,16'd1005,16'd3793};
dout[803]={ -16'd689,-16'd2262,16'd4862,16'd4056,-16'd402,-16'd3366,-16'd5689,-16'd3492,16'd1800,-16'd6498,16'd109,16'd696,-16'd3427,16'd2142,16'd7776,-16'd456,-16'd4874,-16'd4400,-16'd3557,16'd5182,16'd2396,-16'd2264,-16'd6360,-16'd1384,-16'd6719,-16'd8278,-16'd626,-16'd4243,16'd3166,-16'd1185,16'd3395,-16'd1525,16'd3241,16'd5291,16'd2258,16'd4164};
dout[804]={ 16'd5335,16'd5386,16'd2096,-16'd2678,-16'd6335,16'd1434,16'd9080,-16'd5942,16'd3082,-16'd7307,-16'd397,16'd938,-16'd3313,16'd430,-16'd3921,-16'd2907,16'd3755,-16'd564,-16'd4532,16'd1123,-16'd6841,16'd1799,16'd1934,-16'd4122,16'd394,-16'd1874,-16'd11449,-16'd6655,-16'd3264,-16'd2909,-16'd2309,-16'd5368,-16'd561,16'd2210,-16'd1570,-16'd7070};
dout[805]={ 16'd1932,16'd364,16'd469,16'd5099,-16'd4501,-16'd2912,-16'd2875,16'd2026,16'd6964,16'd3241,16'd7334,16'd925,-16'd3340,16'd1941,-16'd7509,-16'd2925,-16'd3699,-16'd5971,16'd5114,-16'd554,-16'd4395,16'd6537,16'd5994,-16'd4439,-16'd3721,16'd4851,16'd61,16'd6540,-16'd556,16'd3941,16'd7061,-16'd769,16'd1141,-16'd5488,16'd368,-16'd885};
dout[806]={ -16'd3140,16'd411,-16'd8701,-16'd7897,-16'd1954,-16'd6159,16'd5465,16'd5543,-16'd642,-16'd3276,16'd2285,16'd5810,-16'd1654,16'd2348,16'd3647,-16'd482,-16'd704,-16'd1326,16'd5879,16'd3666,-16'd624,-16'd683,16'd2170,-16'd1389,-16'd4495,16'd4670,-16'd3265,-16'd6025,-16'd4307,16'd663,16'd1662,-16'd553,-16'd2726,16'd3295,-16'd2813,16'd5214};
dout[807]={ -16'd1324,16'd2951,-16'd6762,16'd3452,16'd4435,16'd3830,-16'd3406,16'd4398,-16'd454,16'd1935,16'd3532,16'd3415,16'd6000,-16'd6209,16'd4346,-16'd5335,16'd853,-16'd2801,16'd5563,-16'd3639,-16'd7382,-16'd910,-16'd1906,-16'd1447,16'd7004,-16'd2741,16'd1967,-16'd2655,-16'd5455,-16'd2891,16'd1530,-16'd2196,-16'd1000,16'd206,-16'd3797,-16'd2630};
dout[808]={ -16'd1731,-16'd7887,16'd1481,-16'd6391,16'd6447,16'd5545,16'd3854,-16'd6287,16'd4468,16'd7725,-16'd6024,-16'd3625,16'd2147,16'd4591,16'd5699,-16'd1142,-16'd2670,16'd2289,-16'd7342,-16'd206,16'd1631,16'd461,16'd3670,16'd8326,-16'd5823,16'd3062,16'd1297,16'd1415,-16'd2243,16'd55,16'd6996,-16'd3698,-16'd2851,-16'd2482,16'd4184,16'd8211};
dout[809]={ -16'd4384,-16'd3,16'd4939,16'd5052,-16'd1766,16'd2969,-16'd4157,16'd1453,16'd2256,16'd5213,-16'd4664,16'd2544,16'd5406,-16'd7530,-16'd3090,16'd3081,16'd1468,-16'd1354,-16'd4447,16'd5746,-16'd4525,16'd1654,-16'd6310,-16'd964,-16'd1314,16'd4683,-16'd1362,16'd2143,-16'd6366,16'd684,16'd3828,-16'd2295,-16'd6967,16'd446,-16'd960,16'd4120};
dout[810]={ -16'd1914,16'd5157,-16'd4416,-16'd4960,-16'd9066,-16'd7130,-16'd400,16'd8844,-16'd143,16'd3132,-16'd3104,-16'd3082,-16'd2024,16'd1855,16'd1856,-16'd2971,-16'd1187,-16'd2074,-16'd3163,16'd2700,-16'd1880,16'd4537,-16'd3587,-16'd2899,16'd2337,16'd2219,16'd862,16'd6840,-16'd4042,16'd9154,16'd2253,-16'd4793,-16'd6515,-16'd6810,-16'd1443,-16'd2981};
dout[811]={ 16'd1978,16'd341,-16'd2870,16'd2443,-16'd3624,-16'd6420,16'd1791,16'd605,-16'd5782,-16'd5152,16'd385,16'd7423,16'd5085,-16'd2980,16'd907,16'd3560,16'd3050,-16'd1892,-16'd1020,16'd2154,-16'd8602,-16'd2650,-16'd5929,16'd5402,16'd29,16'd4580,16'd4821,16'd4772,16'd2151,-16'd8166,16'd5602,16'd2973,16'd5157,-16'd2554,-16'd1974,-16'd6294};
dout[812]={ 16'd6427,16'd5796,16'd2999,16'd2361,16'd3489,16'd721,-16'd3485,-16'd818,16'd2815,-16'd10871,16'd3758,-16'd1802,-16'd5767,-16'd3606,16'd2370,16'd8159,16'd7877,-16'd8006,16'd4485,-16'd6445,16'd6089,-16'd6414,-16'd3410,-16'd9228,-16'd7498,16'd4517,-16'd4070,16'd5351,16'd1041,-16'd4913,16'd6905,16'd8474,16'd635,-16'd8231,-16'd571,16'd4031};
dout[813]={ -16'd2470,16'd8872,-16'd5769,16'd6101,16'd662,16'd6728,-16'd3652,-16'd292,16'd3899,16'd5011,16'd8503,16'd4714,-16'd2804,16'd2532,-16'd3578,-16'd989,16'd2721,-16'd5971,-16'd1942,-16'd2060,-16'd4278,-16'd5251,-16'd1188,-16'd8763,16'd4176,16'd439,-16'd11263,16'd46,-16'd7626,-16'd1883,16'd1147,16'd3217,-16'd190,16'd42,-16'd3693,-16'd6381};
dout[814]={ 16'd4428,-16'd2202,16'd4852,-16'd7181,16'd4513,-16'd8321,16'd9236,-16'd1473,-16'd4052,-16'd3907,16'd4771,16'd7220,16'd1090,16'd2028,16'd6648,-16'd3641,16'd893,-16'd8246,16'd2052,16'd9560,-16'd1495,16'd5047,16'd7083,16'd2870,-16'd5910,-16'd6370,-16'd2676,16'd3536,16'd5782,16'd4601,-16'd9718,-16'd2322,16'd144,-16'd6992,-16'd8706,16'd5921};
dout[815]={ 16'd4976,-16'd3389,16'd2265,16'd2166,16'd2027,-16'd5273,16'd6321,16'd6662,-16'd4077,16'd2294,-16'd1620,-16'd2882,-16'd4240,-16'd4247,-16'd5092,16'd202,-16'd995,16'd5041,-16'd8450,-16'd2001,16'd7188,16'd418,16'd4817,16'd3181,16'd4836,-16'd6562,16'd4580,16'd4754,16'd570,16'd5657,16'd4496,-16'd1612,16'd2245,-16'd4378,-16'd442,16'd3364};
dout[816]={ 16'd6031,16'd3961,-16'd6293,-16'd578,16'd3375,16'd3209,-16'd3092,-16'd3760,16'd928,16'd8129,16'd1331,16'd2533,-16'd1386,-16'd5397,-16'd2243,16'd59,-16'd5125,-16'd2956,-16'd6019,16'd5621,-16'd3459,16'd1987,-16'd2072,-16'd2963,16'd77,16'd1679,-16'd4518,-16'd2608,16'd3020,16'd2135,16'd1696,-16'd5079,-16'd1515,-16'd5852,-16'd5559,-16'd5229};
dout[817]={ 16'd2187,16'd1855,-16'd1780,16'd3129,16'd2853,16'd279,-16'd3923,-16'd4480,16'd2530,-16'd4565,-16'd3560,16'd3556,16'd6771,16'd4003,16'd1521,16'd4693,-16'd330,16'd3210,-16'd6546,-16'd6627,-16'd1364,16'd876,16'd1746,16'd5263,16'd1630,-16'd1207,-16'd4577,16'd1806,16'd7817,16'd6291,16'd5782,16'd5666,16'd4545,-16'd542,-16'd745,16'd5611};
dout[818]={ 16'd4614,-16'd3937,16'd3986,16'd2786,16'd1774,16'd3589,16'd937,16'd5,-16'd2024,-16'd2542,-16'd8233,-16'd7442,-16'd4338,16'd722,16'd5669,16'd3048,-16'd3811,16'd1188,-16'd7735,-16'd1345,16'd5958,16'd4504,16'd4925,16'd2775,-16'd4699,16'd115,16'd2868,16'd2112,-16'd3057,16'd4402,-16'd4453,16'd6194,-16'd1046,16'd1506,-16'd7189,-16'd6990};
dout[819]={ -16'd4543,16'd2235,-16'd808,-16'd705,-16'd6216,-16'd6003,-16'd2790,-16'd6907,16'd168,16'd973,-16'd3264,-16'd4858,-16'd1330,16'd5419,16'd7288,16'd4601,16'd1412,-16'd7576,16'd373,-16'd2084,16'd619,16'd5133,-16'd4031,16'd5303,16'd2846,-16'd3269,16'd3856,16'd5978,-16'd7010,-16'd6574,16'd6009,-16'd2512,16'd2398,16'd439,-16'd1740,16'd1524};
dout[820]={ 16'd400,16'd9386,-16'd5311,16'd438,-16'd8035,16'd3902,-16'd1802,16'd3305,-16'd3011,16'd72,16'd8597,-16'd5856,16'd4657,-16'd2037,16'd289,-16'd1509,16'd5613,-16'd3207,-16'd3501,-16'd4530,-16'd1732,16'd612,16'd1923,-16'd4323,-16'd8337,16'd4366,-16'd7163,-16'd1542,16'd3198,16'd9544,16'd297,-16'd214,16'd6117,16'd305,-16'd149,-16'd1978};
dout[821]={ 16'd5918,-16'd2101,16'd524,16'd173,16'd6869,16'd3040,16'd4751,16'd7855,-16'd6625,-16'd8327,-16'd971,16'd109,16'd2075,16'd3452,16'd3497,16'd4041,16'd5263,-16'd8951,-16'd9049,16'd3392,-16'd3531,16'd3073,-16'd1048,-16'd144,-16'd6870,-16'd8043,16'd6679,-16'd443,-16'd4160,16'd5610,16'd703,-16'd4824,16'd7412,-16'd781,16'd1643,16'd3186};
dout[822]={ -16'd5434,16'd7190,-16'd6911,-16'd3960,-16'd5582,16'd4060,16'd2188,16'd5769,16'd1093,-16'd10580,16'd856,16'd5398,-16'd4373,-16'd4060,-16'd1164,16'd6168,-16'd2411,-16'd5210,16'd6903,-16'd2929,-16'd5244,-16'd5807,16'd2964,16'd1779,-16'd8009,16'd6777,-16'd1240,-16'd3452,-16'd3549,-16'd2834,16'd5534,16'd5388,-16'd2082,-16'd7432,16'd6285,-16'd7268};
dout[823]={ -16'd631,-16'd3156,-16'd5547,16'd5299,-16'd801,-16'd4880,16'd5653,16'd7290,16'd1080,-16'd6893,-16'd2958,16'd7251,16'd3847,16'd1714,-16'd3815,16'd6067,16'd4151,-16'd66,16'd7929,-16'd2050,16'd4535,16'd3907,-16'd5784,-16'd1519,16'd412,-16'd5222,-16'd377,-16'd316,16'd2636,16'd2081,16'd518,16'd2106,16'd2147,-16'd5747,-16'd8384,-16'd4696};
dout[824]={ -16'd3052,16'd4365,-16'd4617,16'd1517,-16'd2803,-16'd1157,16'd2616,16'd7880,-16'd2860,-16'd1883,-16'd3711,16'd2547,-16'd4170,16'd3183,-16'd5739,16'd5288,16'd126,-16'd4756,-16'd7579,-16'd95,-16'd5196,-16'd471,16'd2534,16'd1837,16'd2232,-16'd6162,-16'd5440,-16'd2103,16'd767,-16'd2020,-16'd3848,-16'd3146,-16'd4775,-16'd2513,-16'd9375,16'd4139};
dout[825]={ 16'd4398,16'd3050,16'd1674,-16'd6017,-16'd1673,-16'd2249,-16'd700,-16'd2899,16'd891,-16'd5251,16'd858,-16'd1676,-16'd5134,16'd11,16'd4683,16'd5095,-16'd2314,-16'd4946,-16'd4074,-16'd2392,16'd5487,-16'd4475,-16'd5742,-16'd4218,-16'd8004,16'd6302,-16'd5476,-16'd1106,16'd2259,16'd6815,-16'd2340,-16'd4287,-16'd6270,-16'd7551,16'd500,-16'd8614};
dout[826]={ -16'd7030,-16'd2764,16'd5351,-16'd1723,-16'd4602,16'd1276,16'd1005,16'd1627,16'd59,-16'd550,16'd7099,-16'd6778,16'd3695,16'd705,16'd1443,16'd1935,-16'd721,-16'd5463,-16'd1178,16'd68,-16'd5214,16'd2125,-16'd364,16'd6484,16'd5913,-16'd2258,-16'd1883,16'd2830,-16'd3885,16'd6007,-16'd4669,-16'd5157,-16'd4320,-16'd1744,-16'd342,-16'd2290};
dout[827]={ 16'd2549,16'd1235,-16'd2719,16'd4450,-16'd3646,-16'd5716,16'd1893,16'd644,-16'd3533,16'd2668,16'd4894,-16'd5744,16'd2074,16'd3466,16'd2662,-16'd3531,16'd2858,16'd1714,-16'd5754,-16'd747,16'd5039,-16'd5380,16'd7004,-16'd2821,-16'd7604,16'd4619,16'd4067,16'd2206,16'd6057,-16'd3574,16'd2864,-16'd1455,-16'd7369,-16'd2137,-16'd5252,-16'd4500};
dout[828]={ 16'd5825,16'd5727,-16'd3358,16'd1184,-16'd878,-16'd2696,-16'd999,-16'd7547,16'd4732,16'd6181,16'd4619,-16'd1533,16'd2764,16'd3464,16'd5932,-16'd5256,-16'd4657,-16'd7355,-16'd6663,-16'd2903,16'd1699,16'd4471,16'd4152,16'd872,-16'd6047,-16'd2541,-16'd1290,16'd554,-16'd2261,16'd2701,-16'd2035,-16'd637,16'd1719,-16'd5948,16'd4980,-16'd8188};
dout[829]={ 16'd5996,16'd7905,16'd5878,16'd4431,16'd1038,16'd2137,16'd2252,16'd4514,-16'd3041,-16'd3627,16'd5030,16'd4998,-16'd412,-16'd4184,16'd3448,-16'd7307,-16'd5540,-16'd2039,-16'd4547,16'd3289,-16'd3425,-16'd3001,-16'd5692,16'd1097,16'd2003,-16'd1799,-16'd2553,16'd3429,16'd614,16'd6686,-16'd3476,-16'd2732,16'd2892,-16'd3612,16'd5460,-16'd4632};
dout[830]={ -16'd7143,16'd9343,16'd3365,16'd2011,-16'd4081,16'd2807,-16'd6262,16'd1492,16'd819,16'd2542,-16'd2655,-16'd1048,16'd3983,-16'd3037,-16'd7651,-16'd1059,16'd6388,16'd3695,-16'd6098,-16'd7473,16'd1689,-16'd670,-16'd3150,-16'd4874,16'd625,16'd4316,-16'd5635,16'd597,16'd3184,16'd6933,16'd2905,16'd5450,16'd3777,16'd504,-16'd6418,-16'd1193};
dout[831]={ -16'd7299,-16'd5037,-16'd5549,-16'd267,-16'd5453,16'd2137,-16'd6579,16'd7855,-16'd5492,-16'd4041,-16'd496,-16'd5962,16'd2943,16'd1580,-16'd7188,-16'd6975,-16'd2912,16'd1830,-16'd267,-16'd982,-16'd850,16'd1337,-16'd9016,-16'd6073,-16'd3873,-16'd3015,-16'd489,-16'd4854,-16'd3885,-16'd465,16'd702,16'd7294,16'd4044,-16'd2095,-16'd5942,-16'd2648};
dout[832]={ -16'd8604,-16'd2188,-16'd6510,16'd4784,16'd118,-16'd1564,16'd38,-16'd3714,-16'd8429,-16'd5488,16'd5256,16'd7566,16'd481,16'd3596,-16'd4077,-16'd6062,-16'd7259,-16'd1553,16'd2903,16'd252,-16'd1833,-16'd5568,-16'd293,-16'd2447,-16'd8309,-16'd5855,16'd3791,16'd1031,16'd6814,16'd2142,16'd802,16'd5959,-16'd7001,-16'd5942,16'd4273,-16'd2463};
dout[833]={ -16'd7806,-16'd2470,-16'd5925,-16'd1864,16'd5355,16'd7030,16'd4916,-16'd3536,16'd1254,-16'd762,16'd10025,16'd650,-16'd7091,-16'd1071,16'd3632,-16'd1097,-16'd2648,-16'd540,-16'd1083,-16'd1692,-16'd6733,16'd882,16'd2941,-16'd7404,-16'd5278,-16'd1860,-16'd10085,16'd2238,-16'd3351,16'd2847,16'd9477,16'd1385,16'd2834,-16'd4454,16'd6565,16'd5022};
dout[834]={ -16'd4162,-16'd2513,-16'd2562,-16'd5694,-16'd3493,-16'd6163,16'd7196,16'd1063,16'd1989,16'd10096,-16'd1912,-16'd1516,16'd4680,-16'd1606,16'd1748,-16'd1231,-16'd5007,-16'd1192,-16'd8866,16'd6687,-16'd5080,-16'd1653,-16'd1927,16'd598,16'd2080,16'd540,16'd3745,-16'd5673,16'd898,-16'd373,16'd6089,16'd427,16'd118,16'd2541,16'd4830,16'd1872};
dout[835]={ -16'd395,16'd5729,-16'd7820,16'd4473,-16'd3582,16'd2627,-16'd4921,16'd5127,16'd1181,16'd9442,-16'd5232,-16'd290,-16'd2751,-16'd1560,-16'd2862,16'd2362,16'd435,-16'd2314,-16'd9021,-16'd6031,16'd4860,16'd3685,16'd3407,-16'd7254,-16'd3841,16'd3299,-16'd2255,-16'd1494,16'd5120,-16'd3390,-16'd4426,-16'd2099,16'd324,16'd1314,16'd6655,16'd6009};
dout[836]={ 16'd1567,16'd2527,-16'd6638,-16'd4451,16'd69,-16'd4724,-16'd4269,16'd2909,16'd3805,16'd312,-16'd2598,-16'd9507,16'd4508,16'd5141,-16'd102,-16'd606,-16'd5086,-16'd3502,16'd5310,-16'd6279,16'd3998,16'd4086,16'd5842,16'd4466,16'd2670,16'd6154,16'd6070,-16'd1393,-16'd2933,-16'd2557,16'd293,-16'd7686,-16'd1153,16'd2752,16'd3784,-16'd5756};
dout[837]={ -16'd3706,16'd4232,-16'd3794,16'd6207,-16'd5046,16'd2381,16'd236,16'd3146,16'd675,-16'd4929,16'd1124,-16'd6779,-16'd8405,16'd2456,16'd3263,-16'd5489,16'd917,16'd1601,-16'd4076,16'd5512,16'd1456,-16'd7205,16'd4217,-16'd569,16'd4820,16'd4761,-16'd6712,16'd7121,-16'd3609,16'd2917,-16'd2810,-16'd2767,16'd1746,-16'd7732,16'd1192,16'd114};
dout[838]={ 16'd24,16'd9375,-16'd1158,-16'd3380,-16'd3171,16'd809,-16'd3031,16'd268,16'd2243,-16'd7951,-16'd2305,16'd5170,16'd713,-16'd7634,-16'd6314,-16'd4673,16'd1505,-16'd213,-16'd4725,16'd461,16'd3729,16'd3895,-16'd7351,16'd2358,16'd4952,-16'd6051,16'd2181,16'd5131,-16'd6844,-16'd4642,-16'd7248,-16'd5808,16'd46,16'd4628,16'd7097,16'd3194};
dout[839]={ -16'd2011,16'd412,16'd7375,16'd6609,16'd3994,16'd917,16'd3111,16'd176,16'd2790,-16'd3019,16'd6248,16'd1989,16'd1634,-16'd9820,-16'd6524,-16'd87,-16'd4557,-16'd7981,-16'd3188,16'd3428,-16'd5487,16'd636,16'd6905,-16'd550,16'd4306,-16'd6299,16'd6093,16'd4578,16'd1023,-16'd195,-16'd7692,16'd2702,-16'd194,16'd5726,-16'd1267,16'd1065};
dout[840]={ -16'd1331,-16'd964,16'd853,-16'd7687,-16'd3502,16'd719,16'd6740,16'd10727,-16'd8922,-16'd6866,-16'd423,-16'd1814,-16'd1711,-16'd3308,16'd7543,-16'd1478,-16'd3921,-16'd1160,-16'd7639,-16'd4176,-16'd2963,16'd3182,-16'd1540,16'd791,-16'd5349,-16'd4523,16'd3583,16'd699,16'd5758,16'd3160,-16'd11735,-16'd61,16'd2134,16'd1059,-16'd5256,-16'd3107};
dout[841]={ -16'd6154,-16'd1388,-16'd2497,-16'd3242,16'd5763,16'd9305,16'd1184,16'd3415,16'd4187,-16'd1196,-16'd4617,-16'd4691,-16'd5181,-16'd6548,16'd248,-16'd7421,-16'd7323,16'd4093,-16'd2669,-16'd4413,16'd6985,-16'd3743,-16'd695,16'd5547,16'd3532,-16'd7966,16'd877,-16'd1028,-16'd1218,16'd928,-16'd4443,-16'd1172,16'd5644,-16'd823,-16'd1677,16'd2149};
dout[842]={ -16'd4075,-16'd2763,-16'd4094,16'd4130,-16'd5633,16'd6711,16'd4577,-16'd2555,-16'd1692,-16'd6441,16'd2540,16'd5199,-16'd5621,-16'd1477,-16'd4536,16'd667,16'd5468,-16'd1304,16'd3863,-16'd2703,-16'd6273,-16'd8970,-16'd6639,-16'd3620,-16'd6597,16'd6973,-16'd4497,16'd7768,-16'd2386,16'd752,-16'd6362,16'd5730,16'd462,-16'd775,16'd3252,-16'd4295};
dout[843]={ -16'd6287,-16'd2488,16'd4690,16'd3498,-16'd7017,-16'd1506,16'd1398,-16'd167,-16'd1027,16'd2019,-16'd92,16'd3858,-16'd8723,16'd4345,16'd855,-16'd4156,-16'd3202,-16'd2495,16'd3607,-16'd6884,16'd1386,16'd3536,16'd3259,16'd3854,16'd1273,-16'd641,16'd1450,16'd2465,-16'd3790,16'd4165,-16'd5064,-16'd1580,16'd5963,-16'd8760,-16'd4044,16'd2816};
dout[844]={ 16'd3290,-16'd1898,-16'd2026,16'd518,-16'd7483,16'd3295,16'd3550,16'd92,16'd2615,16'd9075,16'd819,-16'd5799,-16'd4581,16'd3634,16'd1967,16'd7537,-16'd408,-16'd661,16'd3325,16'd2369,16'd6461,16'd6028,16'd3413,-16'd3371,16'd3969,16'd1964,-16'd6075,-16'd900,-16'd888,16'd1575,-16'd3668,16'd5896,-16'd2678,-16'd8398,16'd2470,-16'd645};
dout[845]={ -16'd788,16'd828,-16'd5313,16'd1080,-16'd2190,-16'd1858,16'd3830,-16'd75,16'd1471,16'd9347,16'd6046,-16'd5182,-16'd8416,16'd480,16'd6708,16'd4160,-16'd7187,16'd3383,16'd805,-16'd2065,-16'd223,-16'd6643,16'd2392,16'd810,-16'd7698,-16'd5652,-16'd8502,-16'd6021,-16'd1386,16'd1146,16'd2138,16'd1161,16'd2134,-16'd3678,-16'd4599,16'd350};
dout[846]={ 16'd2401,-16'd1283,16'd1941,16'd4866,16'd1000,-16'd2487,-16'd1247,-16'd7801,16'd2471,-16'd1645,-16'd2442,16'd3733,16'd6117,-16'd2079,-16'd6077,16'd5538,-16'd7658,-16'd3244,16'd4957,16'd365,-16'd5680,16'd3910,-16'd1758,-16'd7382,-16'd8594,-16'd7147,16'd143,16'd6117,-16'd3272,16'd6529,-16'd1960,16'd183,16'd875,16'd4194,16'd5668,16'd5916};
dout[847]={ 16'd2778,16'd2055,16'd4624,16'd1484,-16'd5300,16'd3423,16'd4471,-16'd2280,-16'd1247,16'd2346,16'd3241,16'd1861,-16'd4310,-16'd6155,16'd533,-16'd1585,-16'd2753,16'd6656,16'd5195,16'd7203,16'd1819,16'd4469,-16'd5335,16'd7362,-16'd1727,-16'd5427,16'd2100,16'd5449,-16'd5688,-16'd6167,16'd5765,-16'd4437,-16'd5836,16'd4531,-16'd1665,16'd709};
dout[848]={ 16'd2563,-16'd346,-16'd4805,-16'd6350,-16'd6062,16'd5320,16'd770,-16'd2747,16'd202,-16'd4542,-16'd3387,-16'd3382,16'd3866,16'd4942,-16'd554,-16'd2317,16'd2144,16'd3029,-16'd6243,-16'd1093,-16'd1679,-16'd2640,16'd5227,16'd6592,-16'd307,16'd310,16'd3990,16'd6668,16'd8062,-16'd7069,16'd2616,16'd1591,-16'd1884,16'd1319,-16'd2672,16'd2564};
dout[849]={ 16'd1736,16'd6540,16'd1496,-16'd4032,-16'd3793,16'd5779,-16'd3419,16'd6398,-16'd906,16'd1722,16'd1822,16'd6132,16'd855,-16'd8149,-16'd4927,-16'd3767,16'd7033,16'd5266,16'd2623,16'd7274,-16'd1709,16'd918,16'd163,-16'd839,16'd5429,16'd5099,-16'd7307,-16'd1016,16'd3872,-16'd3057,-16'd5289,-16'd1732,-16'd1346,16'd2664,16'd2544,-16'd6831};
dout[850]={ -16'd4737,16'd10372,-16'd1916,-16'd10572,16'd2950,-16'd4478,16'd2735,-16'd88,-16'd3363,16'd1603,16'd178,16'd768,-16'd4739,16'd6243,-16'd4178,16'd1615,16'd1647,-16'd5457,16'd3377,-16'd184,-16'd3163,16'd613,16'd5119,-16'd6289,-16'd2103,-16'd6535,-16'd7863,-16'd6026,-16'd868,16'd2532,-16'd2150,16'd1367,16'd1907,-16'd9881,16'd1322,16'd1272};
dout[851]={ -16'd298,-16'd7062,16'd6182,-16'd4239,-16'd2904,16'd6735,-16'd3678,16'd246,16'd2022,-16'd2392,16'd1965,-16'd1770,16'd5035,-16'd7476,-16'd2453,-16'd7789,16'd1107,-16'd9598,-16'd6040,-16'd5849,-16'd2432,-16'd8160,16'd3426,16'd6516,16'd2884,-16'd1341,16'd4396,16'd3528,-16'd89,-16'd4224,-16'd2920,-16'd5614,-16'd443,-16'd5621,16'd4699,-16'd4568};
dout[852]={ -16'd2114,16'd4521,-16'd3981,-16'd3715,-16'd2847,16'd5597,16'd6200,-16'd8144,-16'd5941,16'd2080,16'd1565,-16'd389,-16'd6588,-16'd6765,16'd5905,-16'd298,-16'd8953,16'd1818,16'd4904,16'd1349,-16'd492,-16'd11640,-16'd2057,-16'd1831,16'd4789,16'd4329,16'd1697,16'd4931,16'd4616,-16'd5196,16'd263,-16'd5753,16'd3326,16'd2401,16'd2515,16'd3183};
dout[853]={ 16'd11,-16'd2677,-16'd5146,16'd2228,16'd5072,16'd9484,16'd3076,-16'd4864,16'd5816,16'd7765,-16'd5175,16'd3355,-16'd235,16'd8048,-16'd3248,-16'd3287,16'd6406,16'd1784,-16'd2130,16'd4959,-16'd299,-16'd3132,-16'd561,-16'd7677,-16'd2346,-16'd148,-16'd298,-16'd520,16'd5159,-16'd2262,16'd4692,16'd4608,16'd2089,-16'd6880,16'd6432,-16'd5414};
dout[854]={ -16'd7119,-16'd9287,-16'd7577,16'd482,16'd5758,16'd757,16'd733,-16'd4184,-16'd3422,16'd2695,16'd2711,16'd2179,-16'd7349,16'd4996,-16'd5379,16'd567,16'd4112,-16'd390,16'd4978,-16'd27,-16'd6463,16'd552,16'd1324,-16'd2044,-16'd3751,16'd3906,16'd1816,-16'd7572,16'd6573,16'd7187,16'd2317,16'd5152,16'd5732,16'd2026,-16'd185,-16'd570};
dout[855]={ 16'd1890,16'd4798,16'd5314,-16'd1301,-16'd3815,16'd5560,16'd5253,-16'd4347,16'd2480,16'd446,-16'd78,16'd2277,16'd753,16'd3744,-16'd866,16'd4779,16'd5230,-16'd1135,16'd4748,-16'd7991,16'd1107,16'd5709,16'd4064,16'd225,16'd2303,-16'd3787,-16'd8284,16'd4206,16'd5245,-16'd3400,16'd3035,16'd1796,-16'd2736,16'd1952,16'd924,16'd147};
dout[856]={ 16'd7449,-16'd3797,16'd1076,-16'd8284,-16'd1126,16'd1901,-16'd3153,-16'd7616,-16'd3951,16'd3145,16'd504,-16'd9394,16'd6399,16'd5801,-16'd4768,16'd4442,16'd5813,16'd5115,16'd6761,16'd5103,-16'd2717,16'd5001,16'd3754,-16'd1656,-16'd5012,16'd1376,16'd15,-16'd4199,-16'd5595,-16'd1990,-16'd4339,-16'd1937,16'd5195,16'd2285,16'd1724,16'd4139};
dout[857]={ 16'd4818,-16'd7648,16'd1354,16'd5756,16'd3069,16'd3006,16'd3852,-16'd6451,16'd7323,-16'd3852,16'd5422,-16'd6274,-16'd7868,-16'd5823,16'd1836,16'd3556,-16'd5166,16'd4025,16'd4291,16'd786,-16'd662,-16'd1200,-16'd2849,16'd767,-16'd4726,-16'd5155,16'd6667,16'd4589,-16'd4579,16'd6261,16'd4758,16'd1661,16'd6086,-16'd3056,-16'd7763,-16'd333};
dout[858]={ 16'd1442,-16'd924,16'd1445,-16'd4070,16'd3910,16'd3295,16'd1084,16'd4966,-16'd6043,-16'd625,-16'd5005,-16'd3038,16'd2986,-16'd836,-16'd5780,16'd4100,-16'd4201,-16'd4272,-16'd3618,16'd4707,16'd4929,16'd4425,16'd1098,-16'd6217,-16'd1930,16'd7315,-16'd2092,16'd2500,16'd7657,-16'd2823,16'd4237,16'd4060,-16'd8792,-16'd1551,-16'd5803,-16'd910};
dout[859]={ -16'd7516,16'd3815,-16'd4278,-16'd2873,16'd446,-16'd6236,16'd4630,-16'd2399,-16'd4786,-16'd5725,16'd3217,16'd4369,16'd1292,-16'd608,16'd1165,-16'd4002,16'd1890,16'd7469,16'd4423,16'd5843,16'd1833,16'd7267,16'd1168,-16'd5212,16'd2121,-16'd2,16'd1714,-16'd5818,-16'd5536,16'd1794,16'd777,16'd3165,16'd3977,16'd11,-16'd7220,-16'd7262};
dout[860]={ 16'd5161,16'd2298,-16'd2603,-16'd4774,-16'd2408,16'd5331,16'd574,16'd6955,16'd7127,16'd5663,16'd5750,16'd2097,16'd3031,-16'd3201,16'd5386,16'd2749,-16'd9329,-16'd3001,16'd6787,-16'd3019,16'd1786,16'd1047,-16'd3536,16'd6986,16'd5642,-16'd6286,-16'd3053,-16'd5485,16'd104,16'd2004,-16'd11604,16'd1051,16'd3893,-16'd10410,-16'd4077,16'd483};
dout[861]={ 16'd4264,-16'd5955,16'd1736,-16'd2554,-16'd830,16'd7720,16'd3897,16'd2419,-16'd5975,16'd572,16'd5417,-16'd2394,-16'd1973,16'd4674,16'd7326,-16'd9487,16'd620,-16'd7041,16'd2840,-16'd5571,-16'd5600,-16'd2401,16'd5386,16'd1817,16'd4573,16'd472,16'd2656,-16'd1472,-16'd7263,16'd4758,16'd848,-16'd6707,-16'd1967,-16'd8793,16'd1349,16'd4889};
dout[862]={ 16'd4806,16'd4418,16'd4989,16'd7685,16'd6772,-16'd754,16'd6442,16'd766,16'd1269,16'd4875,16'd772,-16'd3941,16'd610,16'd5961,-16'd4821,16'd421,16'd470,16'd4703,16'd2464,-16'd2843,-16'd1845,-16'd4128,-16'd5527,16'd90,-16'd8151,-16'd6659,-16'd340,-16'd4770,16'd6586,-16'd6335,-16'd5208,16'd1685,-16'd7477,16'd5792,-16'd1072,16'd2398};
dout[863]={ -16'd3046,16'd4611,-16'd5664,16'd4913,-16'd405,-16'd1816,-16'd3705,-16'd7556,-16'd8476,16'd6533,16'd4368,16'd4873,-16'd3710,-16'd6486,16'd7628,-16'd1858,16'd1275,16'd3682,-16'd2543,-16'd4902,16'd4251,-16'd7808,16'd4757,-16'd7397,-16'd330,16'd1290,16'd5529,-16'd6037,16'd5925,16'd1215,16'd7170,16'd143,-16'd7242,16'd5788,-16'd4740,-16'd20};
dout[864]={ -16'd1051,-16'd4361,16'd5459,16'd3739,16'd4074,16'd1148,-16'd221,16'd1164,16'd1489,-16'd387,16'd4017,16'd2658,-16'd4835,16'd6726,-16'd162,16'd2165,16'd1214,16'd7452,-16'd6152,16'd3330,-16'd919,16'd3785,16'd183,-16'd5242,16'd2257,16'd5015,-16'd120,16'd3147,-16'd3678,-16'd150,-16'd2738,16'd1719,16'd958,-16'd145,-16'd7536,-16'd6858};
dout[865]={ 16'd1416,-16'd2414,-16'd4040,16'd1064,-16'd1421,-16'd2096,-16'd7473,-16'd2506,-16'd3831,-16'd6354,-16'd4283,16'd2330,-16'd4328,-16'd2527,-16'd5307,-16'd1276,-16'd1488,16'd3851,16'd2372,16'd4585,16'd5600,-16'd98,16'd6151,-16'd7432,-16'd8747,16'd3021,-16'd4251,-16'd423,16'd1982,-16'd2035,16'd5355,16'd6409,16'd6157,-16'd6414,-16'd7210,16'd725};
dout[866]={ 16'd4391,-16'd7666,-16'd7001,-16'd87,16'd1452,16'd4291,-16'd5531,16'd1484,-16'd2,-16'd2559,-16'd4019,-16'd9527,16'd5499,16'd75,-16'd4836,-16'd7836,16'd193,16'd3331,-16'd5399,16'd1939,-16'd387,-16'd1139,-16'd6294,16'd879,-16'd3829,-16'd4543,16'd3787,16'd3231,-16'd6453,-16'd899,16'd665,16'd6293,-16'd4293,-16'd6888,16'd3512,16'd4250};
dout[867]={ -16'd7526,16'd1561,-16'd2904,16'd5107,16'd5138,-16'd6311,-16'd6449,-16'd1696,-16'd1629,16'd7063,-16'd76,-16'd868,16'd746,-16'd6338,-16'd2885,16'd1663,16'd5601,-16'd4838,16'd3226,16'd5668,-16'd196,16'd7628,16'd2234,-16'd3353,16'd1287,16'd250,16'd2388,-16'd3464,-16'd7716,16'd4360,16'd877,16'd2890,-16'd3731,16'd2146,16'd3788,-16'd93};
dout[868]={ -16'd328,-16'd8685,-16'd3791,16'd731,-16'd1697,-16'd6493,16'd1015,16'd6043,16'd2457,16'd1458,-16'd7227,16'd4911,16'd1094,-16'd8246,16'd5476,16'd3221,16'd6953,16'd4267,16'd6895,16'd3836,16'd381,-16'd5937,-16'd1342,16'd3727,-16'd5913,16'd2783,16'd6036,16'd6759,-16'd2315,-16'd5151,16'd3013,16'd5581,-16'd1183,-16'd3098,16'd1049,16'd3832};
dout[869]={ 16'd4078,16'd2835,-16'd1082,16'd1539,-16'd5619,16'd2109,-16'd3918,16'd7000,-16'd991,-16'd3435,16'd5645,16'd3198,-16'd3729,-16'd2768,16'd7437,-16'd2874,-16'd915,16'd7588,16'd6277,-16'd5919,16'd5123,-16'd4099,16'd5633,-16'd3965,16'd1695,-16'd958,16'd4259,16'd323,-16'd4141,16'd230,-16'd1899,16'd1465,16'd1871,16'd619,-16'd4221,16'd4946};
dout[870]={ -16'd669,-16'd5103,16'd4420,-16'd4823,-16'd7688,16'd1430,16'd8301,-16'd2511,16'd2458,16'd1532,-16'd5106,16'd2541,-16'd2557,16'd3946,16'd6038,-16'd5862,-16'd7604,-16'd820,16'd3354,16'd1972,16'd732,16'd5147,-16'd3679,16'd7369,-16'd5895,16'd627,16'd7654,16'd854,-16'd5245,16'd4364,16'd1641,16'd4809,16'd2139,-16'd1068,-16'd4621,-16'd4490};
dout[871]={ 16'd2234,-16'd2036,16'd4725,16'd6508,-16'd6912,16'd1671,-16'd2243,-16'd2355,16'd4424,-16'd3084,-16'd6159,-16'd2770,-16'd5710,16'd2826,16'd3884,16'd1676,-16'd1357,-16'd710,16'd4206,-16'd4775,-16'd5192,-16'd4303,16'd2734,16'd6608,-16'd3633,-16'd4418,-16'd48,16'd3561,-16'd8730,16'd4664,16'd57,-16'd957,-16'd1071,-16'd3684,16'd368,-16'd5771};
dout[872]={ -16'd2963,-16'd5472,-16'd7116,16'd3019,-16'd993,16'd2490,-16'd1751,16'd1002,-16'd1271,16'd6351,-16'd1483,-16'd7509,16'd5166,-16'd4715,16'd7565,-16'd2176,-16'd5698,-16'd3016,16'd1179,-16'd4737,16'd786,-16'd7873,-16'd4640,16'd4516,-16'd3353,16'd3567,-16'd4560,16'd6937,16'd1309,16'd215,16'd1785,-16'd5745,16'd893,-16'd3865,-16'd6911,16'd5606};
dout[873]={ 16'd1567,-16'd9446,16'd6765,16'd2583,16'd6714,16'd2333,-16'd127,16'd4107,-16'd4586,16'd6861,16'd6460,-16'd5654,-16'd4388,16'd2560,-16'd1559,16'd4890,-16'd2105,-16'd8074,-16'd5726,16'd3379,16'd198,-16'd5403,-16'd4306,16'd101,-16'd3210,-16'd1140,16'd483,16'd755,-16'd5951,-16'd4756,-16'd8525,-16'd4345,16'd5613,-16'd723,-16'd6487,-16'd7293};
dout[874]={ -16'd2242,16'd1135,16'd7812,-16'd3460,-16'd4573,16'd7912,-16'd5838,-16'd2182,-16'd748,16'd2778,16'd4750,-16'd6329,-16'd6047,-16'd6733,16'd5813,16'd533,-16'd5577,-16'd1804,16'd4282,16'd6082,16'd3287,16'd297,16'd5114,16'd2303,-16'd3486,-16'd2636,-16'd4534,16'd3033,-16'd2538,16'd8934,16'd5430,16'd5927,16'd4442,16'd2477,16'd1290,16'd2241};
dout[875]={ 16'd3226,-16'd6136,-16'd3094,16'd6584,16'd3461,-16'd3349,16'd3434,-16'd3549,16'd365,-16'd6166,16'd2479,-16'd3008,16'd3957,-16'd5811,16'd3053,-16'd6610,-16'd2135,-16'd5144,-16'd4451,16'd6065,-16'd7231,-16'd5799,-16'd413,-16'd8884,16'd1385,16'd2259,-16'd4634,16'd2439,-16'd1897,16'd2933,-16'd345,16'd2454,16'd6335,-16'd7135,16'd5391,16'd5333};
dout[876]={ 16'd3596,16'd4053,16'd7472,-16'd4756,16'd6058,-16'd1650,-16'd3858,-16'd1531,-16'd5092,-16'd1177,16'd4346,16'd3620,-16'd3267,16'd7784,16'd2572,-16'd3827,-16'd7190,-16'd2328,-16'd3848,16'd3577,-16'd4058,-16'd309,16'd6118,-16'd3219,16'd146,-16'd2603,16'd5395,-16'd4783,-16'd6170,-16'd6600,16'd2148,16'd7251,-16'd6409,16'd7581,16'd3516,-16'd2507};
dout[877]={ -16'd6599,16'd2959,16'd7515,16'd3282,16'd1398,-16'd2292,16'd1788,16'd1461,-16'd7077,-16'd3619,16'd2669,-16'd7425,16'd4143,16'd2478,16'd2642,-16'd7240,-16'd4259,-16'd2556,16'd4901,-16'd1212,-16'd1116,16'd354,16'd2512,16'd5249,-16'd8331,-16'd4144,-16'd2543,-16'd6885,16'd5370,16'd139,16'd4101,16'd6531,-16'd6138,-16'd3462,16'd2108,-16'd1247};
dout[878]={ -16'd579,16'd1327,-16'd6608,16'd5282,16'd934,16'd5265,16'd669,16'd2627,-16'd6969,16'd402,-16'd95,16'd1297,-16'd1316,-16'd3387,16'd4791,-16'd2168,16'd868,16'd1795,16'd1345,16'd581,16'd4870,16'd2195,-16'd1502,16'd4135,-16'd6528,16'd3703,16'd1963,16'd2988,16'd2536,-16'd156,-16'd8258,16'd3937,16'd3497,16'd5528,16'd4802,-16'd3873};
dout[879]={ -16'd5418,-16'd3387,-16'd7125,16'd3329,16'd5355,-16'd3441,16'd4322,16'd2579,-16'd1247,-16'd149,16'd1735,-16'd5026,16'd6184,-16'd2929,-16'd4264,-16'd4747,16'd4123,16'd4680,16'd1106,-16'd3825,16'd550,16'd6245,16'd4695,16'd4728,-16'd4861,16'd3600,16'd4477,16'd4557,16'd4923,16'd4978,-16'd1781,16'd2134,-16'd4793,16'd3731,-16'd1239,16'd5672};
dout[880]={ -16'd4875,16'd7562,16'd6357,-16'd9577,-16'd5054,16'd5102,-16'd1306,16'd3555,16'd6064,16'd9541,16'd453,-16'd2438,-16'd2248,16'd5217,16'd6631,16'd3921,16'd726,-16'd6049,-16'd6281,-16'd2237,-16'd6847,-16'd1316,-16'd3154,-16'd1803,16'd5199,16'd3716,16'd2481,16'd7060,-16'd8312,-16'd356,16'd1881,16'd749,-16'd8346,16'd3592,-16'd8512,16'd2395};
dout[881]={ 16'd7244,-16'd6269,16'd4061,-16'd7152,-16'd5050,16'd2591,-16'd4234,-16'd4324,16'd7819,-16'd5678,16'd353,-16'd1818,16'd804,-16'd1194,16'd804,-16'd10990,-16'd4918,-16'd5214,16'd1590,-16'd4127,16'd3253,-16'd9004,16'd3616,16'd5739,16'd3707,-16'd1511,-16'd1596,16'd7734,16'd5407,-16'd742,16'd1994,-16'd6765,16'd2178,-16'd3096,-16'd6223,-16'd5358};
dout[882]={ 16'd3254,-16'd3345,-16'd7258,-16'd6659,16'd1305,16'd2129,16'd2664,-16'd400,16'd6093,16'd8513,-16'd5841,16'd3419,-16'd1778,-16'd851,16'd4533,-16'd9048,-16'd4256,16'd131,-16'd4770,-16'd10371,-16'd289,-16'd46,16'd2946,16'd3563,16'd4220,-16'd4228,-16'd1271,16'd733,-16'd580,-16'd84,16'd3299,-16'd6220,16'd3473,-16'd6712,-16'd7124,16'd3657};
dout[883]={ -16'd2815,16'd3440,-16'd3970,-16'd7177,16'd2690,16'd8220,-16'd6004,-16'd4516,16'd5264,16'd1109,-16'd1245,-16'd3590,-16'd466,-16'd1404,-16'd372,16'd2838,16'd4404,-16'd2675,16'd6542,-16'd8200,16'd77,-16'd5430,16'd325,16'd6747,-16'd3900,16'd4598,-16'd5705,16'd1288,-16'd6309,16'd5986,-16'd1633,-16'd2493,-16'd1760,-16'd8042,16'd1723,-16'd2410};
dout[884]={ -16'd2631,16'd817,16'd4601,-16'd6347,-16'd6937,-16'd591,-16'd2851,-16'd1804,-16'd3640,-16'd841,16'd4145,-16'd5811,16'd2719,-16'd2272,16'd5959,16'd2258,16'd4680,-16'd4196,16'd5584,16'd1318,-16'd847,16'd968,-16'd2942,16'd5058,-16'd1232,-16'd5381,16'd3080,-16'd6694,16'd310,-16'd1813,-16'd904,-16'd5312,-16'd3084,16'd3666,-16'd4483,16'd711};
dout[885]={ -16'd893,16'd4020,-16'd859,-16'd5732,-16'd148,16'd6826,-16'd7851,-16'd6119,-16'd3254,-16'd523,-16'd2663,16'd2258,-16'd4611,16'd3437,16'd4944,16'd5788,16'd346,-16'd8040,-16'd7786,-16'd598,16'd78,16'd3469,-16'd5575,-16'd3795,-16'd3801,16'd880,16'd4128,-16'd2457,-16'd1593,16'd1353,16'd758,16'd5851,-16'd6197,16'd5259,-16'd14,16'd2084};
dout[886]={ -16'd5582,-16'd7046,16'd2909,16'd4061,-16'd5707,16'd4785,16'd3114,-16'd5549,-16'd6060,16'd7179,-16'd2751,-16'd6201,-16'd4531,-16'd1834,16'd5568,-16'd2352,16'd4149,16'd471,-16'd2363,-16'd4853,16'd6046,-16'd6232,16'd6127,-16'd4895,-16'd6712,-16'd2839,16'd2816,-16'd51,-16'd7437,-16'd5852,16'd117,16'd4771,-16'd3895,16'd1905,-16'd2264,-16'd3088};
dout[887]={ -16'd7079,-16'd5501,16'd7005,16'd7439,-16'd1265,-16'd4397,-16'd4824,16'd5366,-16'd4548,-16'd810,-16'd4593,16'd5895,-16'd6763,-16'd531,16'd6051,16'd2433,16'd3368,16'd2860,-16'd3524,16'd6143,-16'd6467,-16'd1395,-16'd2743,-16'd6943,-16'd289,-16'd2268,-16'd353,16'd308,-16'd5060,16'd414,-16'd6409,-16'd6033,-16'd4133,-16'd4394,-16'd6559,16'd2890};
dout[888]={ -16'd222,-16'd3473,-16'd3998,16'd4665,16'd419,16'd2227,-16'd3917,16'd1196,-16'd7956,16'd7042,16'd5371,-16'd3807,-16'd2333,-16'd2859,-16'd6530,16'd4055,16'd3614,-16'd3095,16'd994,16'd6639,-16'd6040,16'd5639,-16'd2277,16'd3428,-16'd8242,-16'd6402,16'd3487,-16'd1594,16'd4750,16'd5743,16'd1856,-16'd6029,16'd2598,16'd2078,-16'd3443,-16'd2302};
dout[889]={ 16'd1487,-16'd8648,16'd3189,16'd2588,16'd2558,-16'd4338,16'd3086,16'd606,-16'd5031,16'd7119,16'd2937,16'd1266,16'd677,16'd5266,16'd1008,-16'd3632,-16'd6574,-16'd4056,16'd4704,-16'd2199,16'd7001,16'd2596,-16'd4602,-16'd5342,-16'd7299,16'd4670,16'd1396,16'd3238,-16'd3766,-16'd3717,16'd519,-16'd2865,-16'd2374,-16'd5103,16'd1778,-16'd1502};
dout[890]={ -16'd54,16'd983,16'd1402,16'd340,-16'd472,16'd5104,16'd3926,-16'd4733,16'd5462,-16'd1593,16'd2888,16'd181,16'd7811,-16'd7023,-16'd2605,16'd2281,16'd5198,-16'd3421,-16'd6848,16'd3358,16'd4438,-16'd8299,16'd6296,16'd3750,-16'd54,16'd3325,16'd1806,16'd8167,16'd5497,16'd4312,16'd2585,16'd1513,-16'd2441,-16'd6745,16'd1672,16'd2820};
dout[891]={ 16'd3029,-16'd3795,-16'd6329,-16'd6073,16'd3368,16'd8008,16'd307,-16'd9841,-16'd6671,16'd688,-16'd1128,-16'd3808,16'd1889,-16'd4327,16'd5723,-16'd5734,16'd2508,16'd3102,-16'd6289,-16'd3831,-16'd4465,-16'd13163,16'd2739,16'd6638,16'd7673,16'd5521,16'd5961,-16'd2702,-16'd7651,16'd5304,-16'd6860,-16'd362,16'd130,-16'd2330,-16'd9674,-16'd2707};
dout[892]={ -16'd852,16'd4199,16'd1692,-16'd9378,-16'd8175,-16'd1051,16'd5504,-16'd3469,16'd2701,16'd5530,-16'd4901,-16'd2891,16'd3732,-16'd1436,-16'd6942,-16'd8554,16'd5465,16'd3652,-16'd4539,-16'd6069,-16'd1855,-16'd13162,-16'd489,16'd6722,16'd4240,16'd5305,-16'd1072,-16'd2599,-16'd2361,16'd684,-16'd4579,-16'd7728,-16'd3001,16'd4781,16'd5289,16'd2916};
dout[893]={ -16'd1683,-16'd3790,16'd1117,16'd2735,16'd2797,-16'd1933,-16'd9397,-16'd6257,16'd4267,-16'd5198,-16'd2218,-16'd6934,16'd5371,16'd6363,16'd4208,-16'd3992,16'd4375,16'd6239,16'd3870,-16'd96,16'd3812,-16'd2787,-16'd7238,16'd7566,-16'd700,-16'd5306,-16'd363,-16'd9926,16'd3,16'd9113,-16'd5135,16'd6136,16'd2050,-16'd619,-16'd1273,-16'd2769};
dout[894]={ 16'd3276,-16'd5349,16'd1852,16'd2565,-16'd96,16'd4793,-16'd334,16'd5410,16'd5161,-16'd2739,16'd4924,-16'd7368,-16'd7568,16'd3280,-16'd550,16'd4603,16'd3659,-16'd1997,-16'd1446,-16'd6864,-16'd4488,-16'd2624,16'd5422,-16'd4354,16'd7390,-16'd5103,16'd98,-16'd2044,-16'd4736,16'd4526,-16'd2834,-16'd3576,-16'd3290,16'd999,16'd2876,16'd3535};
dout[895]={ -16'd7207,-16'd2466,-16'd4445,-16'd3911,-16'd927,-16'd4245,16'd4589,-16'd6712,-16'd7487,16'd2944,16'd2281,16'd4850,-16'd1122,-16'd154,16'd605,-16'd4577,16'd3151,16'd5031,-16'd1576,16'd5856,-16'd1317,16'd4041,16'd6918,16'd2665,16'd3914,-16'd2750,16'd2675,-16'd4484,16'd644,16'd1351,16'd5576,-16'd7256,-16'd404,-16'd1186,16'd1186,16'd4586};
dout[896]={ -16'd3553,16'd5828,16'd1924,16'd670,-16'd4751,16'd6998,16'd6012,-16'd4136,-16'd5106,16'd6239,16'd3697,16'd4442,16'd6189,16'd4106,16'd705,16'd1319,-16'd786,16'd4938,16'd6868,16'd1355,-16'd51,16'd4247,16'd5551,16'd7967,-16'd5491,16'd5743,16'd2380,16'd5632,-16'd6059,16'd6085,-16'd313,-16'd27,-16'd2692,16'd855,-16'd1000,-16'd3466};
dout[897]={ -16'd6387,-16'd1478,16'd6143,16'd2584,-16'd649,16'd4501,-16'd3435,16'd2153,-16'd1037,16'd1798,-16'd2931,-16'd4931,16'd3171,16'd289,16'd1948,16'd6423,16'd4776,16'd2770,16'd3009,16'd5058,16'd6153,16'd6148,16'd4570,-16'd3035,-16'd3528,16'd3382,-16'd1752,16'd2168,16'd71,-16'd4388,-16'd3174,16'd1147,-16'd5801,16'd4259,16'd1736,16'd1115};
dout[898]={ 16'd108,16'd2608,-16'd364,16'd2180,16'd5964,16'd3898,-16'd838,16'd6621,-16'd6397,-16'd5401,-16'd547,16'd4308,16'd2164,-16'd5233,-16'd3049,16'd4909,16'd2119,16'd6144,16'd5172,16'd1598,-16'd6755,16'd1376,-16'd3352,-16'd570,-16'd4304,16'd3596,16'd2971,-16'd6537,16'd3980,-16'd7268,-16'd2283,16'd2039,16'd6105,-16'd2150,16'd966,-16'd706};
dout[899]={ 16'd6429,-16'd4313,-16'd1408,16'd4747,16'd2325,-16'd4282,16'd8781,16'd6908,16'd4576,16'd3410,-16'd1981,16'd5047,16'd1142,16'd3066,-16'd6019,16'd6649,-16'd1132,16'd431,16'd5860,16'd5292,16'd4339,16'd734,16'd5708,16'd3930,16'd6491,16'd3203,-16'd3581,16'd3886,16'd821,16'd1461,-16'd6220,16'd859,-16'd1716,-16'd848,16'd5169,-16'd795};
dout[900]={ 16'd1788,16'd3540,-16'd6100,16'd4502,-16'd2259,16'd4437,16'd2308,16'd4317,-16'd282,-16'd5811,16'd2462,-16'd7677,16'd2287,-16'd208,-16'd375,-16'd1146,-16'd1231,-16'd3557,-16'd5017,-16'd35,16'd7752,16'd6079,-16'd3426,-16'd2022,16'd5554,-16'd2758,16'd1991,16'd4823,16'd10057,16'd3288,16'd2853,16'd4613,16'd6799,16'd3114,-16'd3662,16'd6119};
dout[901]={ -16'd4832,16'd7535,-16'd5812,16'd726,16'd2111,16'd2582,-16'd9067,16'd5767,16'd3843,-16'd6195,-16'd7530,-16'd2533,-16'd4812,16'd4898,16'd667,16'd5551,-16'd4519,-16'd4849,16'd4223,16'd7503,16'd6358,-16'd6235,16'd3688,-16'd782,16'd5088,16'd2535,16'd2601,-16'd1912,16'd8057,16'd1315,16'd4129,16'd1155,16'd4335,16'd3308,16'd1114,16'd948};
dout[902]={ 16'd4425,16'd1333,-16'd1217,16'd4582,-16'd7792,16'd4021,16'd289,16'd6841,16'd5478,-16'd10226,16'd3228,-16'd1975,16'd1517,16'd7696,16'd3677,16'd3953,-16'd205,-16'd10883,16'd5753,-16'd9029,16'd8017,-16'd483,16'd4414,-16'd5297,-16'd2617,-16'd4819,-16'd10339,-16'd5772,-16'd3580,-16'd2585,-16'd1820,-16'd1385,-16'd3347,16'd4135,-16'd4953,16'd3333};
dout[903]={ 16'd5731,16'd3682,16'd4476,-16'd3903,-16'd8523,-16'd5009,-16'd581,-16'd4598,16'd617,-16'd6316,16'd5501,16'd622,-16'd3812,16'd3073,-16'd3536,16'd7973,-16'd7258,-16'd2775,16'd7142,-16'd596,16'd5729,16'd8516,-16'd6570,-16'd14425,16'd4277,16'd7311,16'd2606,-16'd1652,-16'd3253,16'd1739,-16'd4524,-16'd5138,16'd3316,16'd3098,-16'd2258,16'd2868};
dout[904]={ -16'd1225,16'd1452,-16'd2973,16'd5600,16'd2820,-16'd3933,16'd5467,-16'd4458,16'd3371,-16'd9983,16'd1655,16'd5217,-16'd1685,-16'd539,-16'd7206,-16'd3095,16'd5181,-16'd2107,16'd1062,-16'd983,16'd2700,16'd2256,-16'd1877,-16'd11690,-16'd1704,16'd2011,16'd3016,-16'd5915,-16'd3701,-16'd643,16'd822,16'd1713,-16'd7660,16'd2472,-16'd4277,-16'd3118};
dout[905]={ -16'd5993,16'd5811,16'd1523,-16'd844,16'd4358,16'd4506,-16'd2375,-16'd3723,-16'd6891,16'd1759,16'd1130,16'd101,16'd2813,16'd2409,16'd1070,-16'd5950,16'd281,-16'd3131,-16'd1787,16'd8949,16'd4448,16'd5333,-16'd2558,-16'd4649,-16'd1641,16'd2098,-16'd3354,-16'd2526,16'd684,-16'd5453,-16'd3958,16'd2627,-16'd4207,-16'd5881,-16'd530,16'd7785};
dout[906]={ -16'd7091,-16'd509,16'd3084,16'd4219,16'd2613,-16'd4686,16'd1655,-16'd3973,-16'd2825,16'd5079,16'd1133,-16'd6466,16'd6921,16'd1111,-16'd3923,-16'd6883,-16'd8609,16'd1358,16'd9220,16'd1003,16'd246,-16'd281,16'd3555,-16'd5338,16'd4193,-16'd8086,16'd5240,16'd4719,-16'd5692,-16'd3691,16'd1467,16'd198,-16'd1027,16'd5720,-16'd2743,16'd8156};
dout[907]={ -16'd4908,16'd6894,16'd3629,-16'd2925,16'd433,-16'd1271,-16'd6802,16'd2588,-16'd6267,16'd5624,16'd4488,16'd7372,16'd7006,-16'd2376,-16'd1248,16'd4457,16'd3095,-16'd1412,16'd6221,-16'd4564,16'd2839,-16'd1654,16'd2070,16'd1555,16'd5993,-16'd3374,-16'd6071,-16'd364,16'd1026,-16'd4645,16'd6010,-16'd805,-16'd4269,16'd6152,-16'd6424,-16'd5602};
dout[908]={ -16'd3879,-16'd1410,-16'd1851,16'd1175,-16'd4064,-16'd3675,-16'd6675,-16'd1650,16'd4106,16'd2597,-16'd580,16'd1142,-16'd558,16'd2725,-16'd1840,16'd1582,16'd2771,16'd6089,16'd2629,16'd1547,-16'd2881,-16'd612,16'd288,16'd3951,16'd8582,16'd4710,16'd3558,16'd3963,-16'd6946,16'd964,16'd2158,16'd4057,-16'd4009,-16'd5313,-16'd6274,-16'd3400};
dout[909]={ 16'd936,16'd866,-16'd606,-16'd681,16'd276,16'd114,16'd6345,16'd5053,16'd5926,16'd3153,-16'd5097,16'd5033,16'd8302,16'd132,-16'd3678,-16'd3453,16'd3378,-16'd8338,16'd2719,-16'd5853,-16'd4309,-16'd3855,16'd6078,16'd1456,16'd1316,-16'd5017,16'd2333,-16'd3555,-16'd3101,16'd9125,16'd3219,16'd3876,-16'd1658,16'd6070,-16'd4169,16'd559};
dout[910]={ -16'd2630,-16'd4923,16'd2504,-16'd1569,-16'd817,-16'd3060,-16'd6253,-16'd2349,-16'd2973,16'd3376,16'd9556,-16'd2124,16'd6549,16'd3668,-16'd717,-16'd1996,-16'd4771,16'd2542,16'd3674,16'd384,-16'd845,16'd5796,-16'd7462,-16'd876,-16'd527,-16'd405,-16'd7826,-16'd4162,-16'd1139,-16'd5523,-16'd4576,-16'd181,-16'd776,16'd365,-16'd6477,-16'd3398};
dout[911]={ 16'd3338,-16'd3144,-16'd4558,-16'd6752,16'd2636,-16'd8607,16'd1608,16'd6497,16'd857,-16'd3455,-16'd5523,16'd3642,-16'd5500,-16'd7528,16'd4934,16'd6637,-16'd647,-16'd10909,-16'd3911,-16'd3606,-16'd5933,16'd6426,-16'd3071,-16'd2507,-16'd5750,16'd1832,-16'd1524,16'd3850,16'd2032,16'd3910,16'd1001,16'd5409,-16'd7743,-16'd3363,-16'd5579,-16'd4588};
dout[912]={ -16'd4892,-16'd7298,-16'd6095,16'd4829,-16'd1149,16'd3734,16'd7958,16'd3795,16'd687,-16'd2242,-16'd6124,16'd7412,-16'd2492,-16'd172,-16'd1775,16'd1302,16'd5366,-16'd6461,16'd2512,16'd5100,-16'd1399,-16'd2001,16'd10378,-16'd7111,16'd63,16'd5542,-16'd780,-16'd469,-16'd3471,16'd2057,-16'd5613,-16'd4167,16'd1324,16'd4208,16'd219,16'd1156};
dout[913]={ -16'd897,16'd6713,16'd3276,-16'd2136,-16'd5035,-16'd1426,-16'd2803,16'd3572,16'd2254,-16'd6638,-16'd6278,16'd7060,-16'd4085,-16'd2052,16'd535,-16'd3514,-16'd5667,-16'd1941,16'd7154,-16'd1803,-16'd1150,16'd306,16'd2218,-16'd3633,16'd5735,-16'd2162,-16'd358,16'd7784,16'd1699,16'd3498,-16'd6886,16'd3604,16'd1694,16'd1875,-16'd8248,16'd4845};
dout[914]={ 16'd6701,16'd6233,-16'd5578,16'd7111,-16'd127,-16'd1371,16'd2083,16'd1085,16'd3098,16'd4031,-16'd586,-16'd607,16'd465,16'd3955,-16'd3111,-16'd114,-16'd7600,16'd124,16'd6480,-16'd4265,-16'd6925,-16'd3448,-16'd10289,-16'd3193,16'd791,-16'd1503,-16'd1083,-16'd5977,-16'd191,-16'd658,-16'd1851,-16'd1495,-16'd5733,-16'd4853,-16'd8215,16'd2000};
dout[915]={ -16'd1109,16'd4077,-16'd6397,16'd1611,-16'd297,-16'd5683,16'd1504,-16'd7534,16'd4000,16'd3476,-16'd3099,16'd1677,16'd2786,16'd6098,-16'd2652,16'd3603,16'd3291,16'd2801,16'd2147,-16'd765,-16'd4746,-16'd1981,-16'd2181,16'd2515,-16'd4279,16'd3262,-16'd788,16'd2088,-16'd388,16'd6602,16'd7386,16'd4048,16'd896,-16'd118,16'd3096,-16'd3942};
dout[916]={ 16'd16,-16'd6122,-16'd7312,-16'd6476,16'd2474,-16'd3211,-16'd1452,16'd4755,16'd5920,-16'd2033,16'd6664,-16'd1211,-16'd5813,-16'd4169,16'd2090,16'd1520,16'd2079,16'd5734,-16'd3506,-16'd3118,-16'd5149,16'd4235,-16'd8338,-16'd1331,16'd911,-16'd4976,16'd1565,-16'd1038,16'd2548,-16'd2033,16'd8512,-16'd1098,16'd3744,16'd5666,-16'd2829,16'd3990};
dout[917]={ -16'd2239,-16'd5097,-16'd4747,-16'd5577,16'd6242,-16'd873,-16'd4351,-16'd7082,-16'd2955,16'd3586,16'd2169,-16'd1013,-16'd3499,-16'd6104,-16'd5043,16'd387,16'd4104,16'd8137,-16'd1586,16'd6225,-16'd2661,-16'd3325,-16'd2153,16'd5352,-16'd1845,16'd2882,16'd2190,16'd4725,-16'd1293,16'd2504,16'd3037,-16'd3239,16'd2760,16'd2551,16'd4989,-16'd5809};
dout[918]={ -16'd6651,16'd144,16'd6129,16'd9068,16'd4104,-16'd8560,16'd1129,16'd4485,-16'd3482,16'd7135,16'd5491,-16'd32,-16'd553,16'd6302,-16'd78,-16'd1904,-16'd8157,-16'd1368,-16'd1765,-16'd514,16'd2845,16'd2074,-16'd6133,16'd5642,-16'd3455,-16'd7506,16'd3941,-16'd820,-16'd1499,-16'd3952,16'd1591,16'd6222,-16'd5115,-16'd1782,-16'd7072,-16'd2862};
dout[919]={ -16'd7393,-16'd4268,16'd159,16'd1224,16'd2064,16'd1897,-16'd6466,16'd3816,-16'd6100,16'd4072,-16'd3949,16'd7195,-16'd2077,-16'd6796,16'd1193,16'd427,16'd134,-16'd2295,16'd2189,-16'd4761,16'd3607,16'd2311,-16'd2170,16'd5331,16'd7229,-16'd6227,16'd1243,16'd6742,-16'd6669,-16'd3526,16'd2962,16'd2613,16'd1659,-16'd4173,16'd6049,16'd2277};
dout[920]={ -16'd2392,-16'd3676,-16'd6320,-16'd5752,-16'd8787,-16'd3453,16'd4581,16'd1451,16'd3437,-16'd7865,16'd3769,-16'd1261,16'd1551,-16'd1643,-16'd5877,16'd3826,-16'd8171,16'd2894,-16'd3466,-16'd4836,16'd2036,-16'd4279,-16'd8862,16'd12221,-16'd2979,-16'd3910,-16'd580,-16'd7425,16'd2101,-16'd7048,16'd7541,-16'd1874,-16'd1004,16'd5515,16'd7315,-16'd6209};
dout[921]={ 16'd3360,16'd1875,-16'd3407,-16'd801,16'd2325,16'd2199,-16'd1331,-16'd4445,-16'd7416,16'd2186,-16'd7506,16'd6453,-16'd8906,-16'd5438,16'd2327,16'd2468,16'd2124,-16'd10542,-16'd2499,16'd7830,-16'd2636,16'd874,16'd2765,-16'd6689,-16'd7255,-16'd3655,16'd1861,16'd820,16'd1773,-16'd576,-16'd829,-16'd782,16'd189,16'd8982,-16'd6007,16'd3086};
dout[922]={ 16'd3358,-16'd4091,-16'd2114,-16'd1921,-16'd1445,-16'd5982,-16'd1592,16'd1051,-16'd8122,-16'd704,-16'd1910,16'd5391,-16'd4258,16'd2971,16'd1282,-16'd1881,16'd1331,-16'd12503,16'd4277,-16'd4019,-16'd1584,16'd3525,16'd899,-16'd820,16'd2187,16'd742,-16'd10063,16'd1439,-16'd822,-16'd5089,-16'd3924,16'd461,-16'd6434,-16'd5402,-16'd3945,-16'd3208};
dout[923]={ -16'd3563,16'd2653,16'd1393,-16'd881,-16'd186,-16'd2047,16'd7340,-16'd1661,16'd1208,16'd4945,16'd1412,-16'd6259,16'd5571,-16'd3562,16'd2524,-16'd1066,16'd4750,16'd1638,16'd1332,-16'd1822,-16'd2819,-16'd866,16'd9478,-16'd2773,-16'd2326,16'd3981,-16'd451,16'd6787,16'd2876,-16'd4570,16'd892,-16'd3126,-16'd7980,16'd9690,16'd6824,16'd4574};
dout[924]={ 16'd8342,16'd5477,-16'd5642,-16'd5622,-16'd828,-16'd4910,-16'd5405,16'd2122,-16'd2859,16'd2820,16'd4191,16'd2956,-16'd6241,16'd9858,16'd587,16'd2650,16'd919,16'd8282,-16'd249,16'd696,-16'd3624,-16'd3319,-16'd5451,-16'd1073,-16'd8942,-16'd1038,-16'd4387,16'd4769,16'd5521,-16'd8435,16'd1566,16'd1290,-16'd3000,16'd1179,-16'd5346,16'd2381};
dout[925]={ 16'd1679,-16'd4519,-16'd7403,16'd531,16'd521,16'd1912,-16'd6952,16'd3613,-16'd2796,16'd478,16'd2307,16'd3137,-16'd7424,-16'd8183,-16'd3443,16'd576,16'd3882,16'd6738,16'd2794,16'd4015,16'd615,16'd4971,-16'd2947,-16'd7260,-16'd4287,16'd6271,16'd3336,16'd3246,-16'd2618,-16'd9296,16'd2827,16'd6487,-16'd3684,16'd1445,16'd388,16'd2481};
dout[926]={ 16'd5846,-16'd5057,16'd1958,-16'd236,-16'd3112,16'd5454,-16'd2129,16'd4277,-16'd7151,-16'd5898,-16'd4589,16'd6465,16'd5013,16'd5162,-16'd10,16'd2204,-16'd3492,16'd8372,-16'd2188,16'd7736,16'd5744,-16'd2260,-16'd4764,16'd2778,16'd3918,16'd4164,-16'd7241,16'd4686,-16'd102,-16'd7809,-16'd4005,-16'd781,-16'd8270,-16'd209,16'd6097,-16'd3752};
dout[927]={ 16'd5579,-16'd638,16'd2796,16'd2348,16'd1261,-16'd4994,-16'd4750,16'd5857,16'd2769,-16'd5939,16'd6249,16'd3269,16'd773,-16'd6028,16'd1072,16'd117,16'd2760,-16'd1030,16'd4106,-16'd4822,16'd5473,-16'd4304,-16'd4439,16'd2571,-16'd2623,-16'd2243,16'd1621,16'd453,-16'd3418,16'd6808,16'd1381,16'd673,-16'd3697,-16'd4421,16'd1060,-16'd2303};
dout[928]={ -16'd7550,-16'd4856,-16'd5083,16'd1106,16'd2955,-16'd11526,-16'd8578,16'd4916,16'd1610,-16'd4281,-16'd6063,-16'd2616,-16'd2329,16'd4757,16'd977,-16'd910,16'd330,16'd3812,-16'd7093,-16'd1016,-16'd4955,-16'd237,-16'd3588,16'd6009,-16'd2361,-16'd3376,16'd1249,16'd782,-16'd7881,-16'd2378,16'd1654,16'd1783,-16'd6368,16'd6593,16'd66,16'd3175};
dout[929]={ 16'd3885,16'd3707,-16'd1067,-16'd2606,16'd3803,16'd4133,16'd3676,-16'd5254,-16'd6454,16'd4735,-16'd7513,-16'd4986,16'd5435,16'd6651,16'd1602,16'd4491,16'd2170,16'd2146,16'd1638,16'd4949,16'd843,16'd7015,-16'd4882,-16'd6464,16'd3221,-16'd4962,16'd454,16'd4488,-16'd4211,16'd5078,16'd3155,16'd2318,-16'd4022,-16'd2097,-16'd4122,16'd438};
dout[930]={ 16'd1341,-16'd687,-16'd2775,16'd598,-16'd5226,-16'd6046,-16'd3374,16'd68,-16'd10796,16'd8148,-16'd1721,16'd3434,16'd2408,16'd545,16'd772,-16'd5190,-16'd1974,-16'd757,-16'd3729,16'd7652,16'd972,-16'd6593,-16'd3339,16'd2953,-16'd5658,16'd5704,-16'd9801,16'd2059,16'd14236,-16'd2195,-16'd187,16'd9046,16'd6776,-16'd3836,16'd130,16'd2586};
dout[931]={ -16'd4276,-16'd6157,-16'd3903,-16'd5187,16'd385,16'd2206,-16'd942,-16'd4231,-16'd1362,16'd254,-16'd3516,-16'd6301,-16'd5441,-16'd1773,-16'd713,16'd4913,-16'd5979,-16'd7513,16'd1390,16'd5122,16'd6105,-16'd2638,16'd4780,-16'd7140,16'd6494,16'd5405,-16'd254,-16'd7147,16'd2701,16'd1913,16'd4415,16'd4136,-16'd2824,16'd3967,16'd275,16'd4997};
dout[932]={ 16'd786,-16'd7301,-16'd3564,-16'd4467,16'd456,-16'd1125,-16'd708,16'd4894,-16'd1192,16'd4735,-16'd9269,16'd1735,16'd1125,16'd4477,16'd1288,-16'd2755,-16'd2417,-16'd1981,16'd1048,16'd3104,-16'd2351,16'd8471,16'd1564,16'd5279,16'd7530,-16'd2773,-16'd8667,-16'd2831,-16'd788,-16'd5505,-16'd5125,-16'd133,16'd5301,-16'd3689,-16'd6407,-16'd9309};
dout[933]={ 16'd31,-16'd7319,16'd1610,-16'd3296,-16'd5119,16'd5947,16'd4758,16'd76,16'd3081,16'd2327,16'd788,-16'd3178,16'd2374,16'd2888,-16'd2860,16'd151,-16'd6010,-16'd2266,-16'd917,-16'd10861,-16'd7374,-16'd3869,-16'd5134,-16'd2134,-16'd8969,-16'd6670,-16'd1030,16'd2449,-16'd5647,-16'd8529,16'd3242,-16'd2369,16'd1423,16'd6333,16'd2119,16'd6410};
dout[934]={ -16'd2666,-16'd2214,16'd1346,-16'd5888,-16'd8182,-16'd804,16'd8121,-16'd416,16'd5873,-16'd4344,16'd2209,-16'd2321,-16'd3625,-16'd30,-16'd5166,16'd7058,-16'd5677,16'd371,16'd3754,-16'd3030,16'd2897,-16'd653,-16'd2,-16'd6225,-16'd7045,16'd4175,-16'd273,-16'd1240,16'd6110,16'd4057,16'd1414,16'd1366,16'd4947,16'd6753,-16'd8251,-16'd5376};
dout[935]={ 16'd6739,-16'd4046,-16'd9215,-16'd2313,16'd4276,-16'd2031,-16'd3227,-16'd6073,16'd7680,-16'd6303,-16'd7052,-16'd1285,-16'd2109,-16'd4961,-16'd607,16'd3388,-16'd2768,16'd7383,-16'd5646,16'd5841,-16'd2297,-16'd2872,16'd4287,16'd4079,-16'd5315,16'd925,16'd7558,16'd4973,16'd7335,16'd4141,-16'd4198,16'd466,-16'd2453,16'd3477,16'd5327,-16'd2345};
dout[936]={ -16'd588,-16'd4260,16'd5742,-16'd666,16'd703,16'd3299,16'd4889,16'd815,16'd2054,16'd7516,16'd4448,16'd2316,16'd4229,-16'd5116,-16'd6220,-16'd5434,16'd759,16'd8251,16'd358,16'd9890,16'd2773,16'd7576,-16'd1942,-16'd1616,-16'd6416,16'd714,16'd4704,-16'd5723,-16'd3482,16'd6080,-16'd4182,-16'd95,-16'd1257,-16'd4730,16'd2975,16'd3781};
dout[937]={ -16'd7794,-16'd3755,-16'd3824,-16'd1413,-16'd1281,16'd4518,16'd5760,-16'd724,-16'd3555,-16'd6319,-16'd1797,16'd5186,16'd2800,16'd2387,16'd262,-16'd2953,16'd4400,-16'd2965,-16'd5261,-16'd5159,16'd2481,-16'd2251,-16'd4481,-16'd4992,16'd5789,16'd3161,16'd6359,16'd3892,-16'd2870,16'd4787,16'd2215,16'd2068,-16'd4882,16'd6127,-16'd8526,-16'd2244};
dout[938]={ 16'd145,-16'd5201,-16'd5481,-16'd5743,-16'd5180,-16'd9688,-16'd5206,-16'd1900,16'd4822,16'd2503,-16'd5985,-16'd4406,16'd3031,16'd792,-16'd6548,-16'd5343,16'd9139,-16'd80,-16'd1626,16'd1800,16'd3138,16'd2292,-16'd164,16'd2016,16'd4201,-16'd6368,16'd6891,16'd2428,16'd5191,-16'd6614,16'd196,16'd1304,-16'd105,16'd5116,-16'd3273,-16'd1585};
dout[939]={ 16'd3612,16'd734,-16'd2023,16'd4679,16'd4672,-16'd1984,-16'd375,-16'd2014,16'd672,-16'd4564,-16'd461,-16'd1004,16'd567,-16'd5801,16'd957,16'd5870,16'd1201,-16'd3024,16'd5652,16'd2445,-16'd5747,16'd1090,-16'd2440,16'd6729,-16'd2220,-16'd3613,-16'd5919,16'd6377,-16'd1038,16'd512,16'd4949,-16'd4060,-16'd2303,16'd3176,16'd2418,-16'd3774};
dout[940]={ 16'd4919,16'd1769,-16'd2445,16'd4636,-16'd6883,-16'd7011,-16'd922,-16'd3596,-16'd3606,16'd3306,16'd2591,16'd1689,16'd6220,16'd2226,16'd2586,16'd4274,16'd3706,-16'd2008,16'd779,-16'd1274,-16'd5091,-16'd5820,16'd288,16'd10204,-16'd852,-16'd1880,16'd6126,16'd1259,16'd8164,-16'd774,16'd8738,-16'd1904,16'd254,-16'd103,-16'd4214,16'd4374};
dout[941]={ -16'd3371,16'd1607,-16'd5165,-16'd5473,16'd2393,-16'd4924,-16'd569,16'd788,-16'd2064,16'd2917,-16'd8682,16'd4973,16'd5361,16'd592,-16'd4281,16'd3304,16'd5936,-16'd5442,16'd3115,16'd3528,-16'd199,-16'd7616,-16'd5662,-16'd4031,16'd3413,-16'd2943,-16'd7847,16'd242,16'd5188,16'd3157,16'd2327,-16'd5509,-16'd155,16'd6133,-16'd337,16'd2922};
dout[942]={ -16'd1952,16'd1388,16'd3194,16'd827,-16'd3682,16'd6557,16'd7064,16'd5290,-16'd4391,16'd4140,-16'd6501,-16'd5429,16'd6948,-16'd2599,16'd5612,-16'd1541,16'd6251,-16'd4221,-16'd2839,-16'd5620,-16'd5156,16'd2331,16'd4580,-16'd2422,16'd5303,-16'd9756,-16'd3351,-16'd6260,-16'd8257,16'd7834,-16'd1832,16'd2553,16'd6848,16'd6862,16'd2297,16'd5212};
dout[943]={ -16'd3701,-16'd906,16'd8220,-16'd507,-16'd1548,16'd2678,-16'd93,16'd6066,16'd335,-16'd692,16'd423,-16'd4951,16'd5594,16'd9048,16'd5509,16'd3784,-16'd602,-16'd5652,16'd6457,16'd467,-16'd5918,-16'd5555,16'd6992,-16'd769,-16'd6737,-16'd4546,-16'd6894,16'd5049,16'd3988,-16'd4043,-16'd6239,-16'd3472,16'd5876,16'd1932,-16'd2356,16'd3618};
dout[944]={ 16'd2090,-16'd4472,-16'd3394,-16'd2070,16'd1301,-16'd4825,-16'd649,16'd4622,-16'd3164,16'd1723,-16'd4510,16'd866,16'd3921,16'd6434,-16'd4847,-16'd4659,-16'd347,16'd2558,-16'd7029,-16'd2365,16'd6356,16'd7089,-16'd2601,-16'd5941,-16'd81,16'd366,-16'd2579,16'd7229,16'd7463,-16'd2490,-16'd7982,-16'd8301,-16'd8153,16'd2963,-16'd7593,-16'd3729};
dout[945]={ -16'd2027,-16'd6108,-16'd4536,-16'd5803,-16'd3649,-16'd1107,16'd5724,-16'd3867,-16'd6891,16'd1539,16'd3860,-16'd2364,16'd5029,-16'd3598,16'd74,-16'd6714,16'd4783,-16'd720,-16'd1247,16'd5403,-16'd4836,-16'd5883,-16'd189,-16'd4835,16'd735,16'd2914,-16'd3015,16'd1596,16'd3328,-16'd4318,16'd8483,16'd3623,16'd1738,16'd6681,16'd4712,-16'd5979};
dout[946]={ 16'd6491,-16'd7071,-16'd4269,16'd1227,-16'd2420,16'd1080,-16'd5955,16'd5125,16'd3728,16'd68,-16'd891,16'd2435,16'd2197,16'd5355,16'd3925,16'd6469,-16'd4192,16'd5690,-16'd5183,-16'd3343,16'd7324,-16'd3293,-16'd93,-16'd777,16'd3138,-16'd4057,16'd5981,-16'd6683,-16'd2370,-16'd6639,-16'd1204,-16'd6866,-16'd7631,16'd5029,-16'd4751,-16'd4441};
dout[947]={ 16'd5212,16'd5884,-16'd7277,16'd2907,16'd4274,16'd4315,-16'd5752,16'd2863,-16'd3304,16'd1860,16'd1374,-16'd6712,16'd5087,16'd4988,-16'd2693,-16'd5606,-16'd6952,16'd5349,16'd854,16'd2064,16'd9686,-16'd3028,-16'd2159,-16'd5187,16'd4409,-16'd3306,-16'd319,16'd4895,16'd780,16'd4763,16'd5193,-16'd758,-16'd3446,16'd1723,16'd3294,16'd7172};
dout[948]={ -16'd4406,16'd1569,16'd3772,-16'd520,-16'd344,-16'd6102,16'd5992,-16'd1426,16'd4118,16'd4890,-16'd3391,16'd3606,16'd4198,-16'd6837,-16'd5282,-16'd1580,16'd700,16'd1291,16'd2153,-16'd1590,-16'd4705,16'd4228,-16'd7850,-16'd6680,16'd6774,-16'd2593,16'd4011,16'd2590,16'd4982,16'd3591,-16'd4869,-16'd6010,-16'd8455,16'd2382,16'd2605,16'd5465};
dout[949]={ -16'd6348,16'd3090,16'd982,16'd1295,16'd5548,16'd272,16'd5187,-16'd868,-16'd4418,-16'd6100,16'd7143,-16'd1754,-16'd249,16'd2863,-16'd6803,16'd6558,-16'd3079,-16'd1245,-16'd7835,-16'd1266,-16'd4278,-16'd4866,-16'd800,-16'd5810,-16'd5476,-16'd3185,-16'd4926,16'd1151,16'd5860,-16'd546,16'd4395,16'd5715,16'd569,16'd3956,-16'd1482,16'd1517};
dout[950]={ 16'd1725,16'd6662,-16'd895,-16'd6722,-16'd2475,16'd2404,-16'd3604,16'd7854,16'd2504,16'd6458,16'd3309,16'd781,16'd3493,16'd6139,-16'd3612,-16'd7504,16'd620,-16'd19,-16'd3970,-16'd59,-16'd4190,16'd2568,-16'd6811,-16'd755,16'd1291,16'd1040,16'd4799,16'd2722,16'd11831,-16'd1797,16'd1193,-16'd5927,16'd2577,-16'd652,16'd6073,-16'd995};
dout[951]={ -16'd4581,16'd892,-16'd2830,-16'd1288,-16'd3329,16'd8476,-16'd1284,-16'd5199,16'd1576,16'd1703,-16'd8462,16'd3332,16'd6065,16'd3631,16'd4219,-16'd8629,-16'd6099,-16'd981,16'd4734,16'd6485,16'd1603,-16'd5706,16'd6190,16'd2767,16'd5791,-16'd1258,-16'd3037,-16'd2330,16'd5335,16'd8181,-16'd2611,-16'd7765,-16'd6330,-16'd1850,-16'd4985,-16'd4693};
dout[952]={ 16'd3476,16'd5812,16'd55,-16'd7794,-16'd1393,-16'd1721,16'd8783,-16'd472,16'd1229,16'd3561,-16'd3813,-16'd4535,16'd1267,-16'd6835,-16'd1139,16'd4356,-16'd8742,16'd515,16'd4976,16'd6695,-16'd1172,-16'd2550,16'd5734,16'd2766,16'd7839,-16'd2194,16'd1544,-16'd11010,-16'd4962,-16'd3771,16'd4667,-16'd7369,-16'd2162,16'd2383,-16'd3587,-16'd4299};
dout[953]={ -16'd7685,-16'd2741,16'd2107,-16'd8298,-16'd531,16'd3725,16'd5340,16'd324,-16'd5341,-16'd555,16'd1797,-16'd1774,16'd3222,-16'd248,-16'd857,16'd7569,-16'd5168,-16'd5953,-16'd289,-16'd4188,16'd5759,-16'd4677,16'd387,16'd7573,16'd2797,16'd4179,16'd3375,-16'd6042,16'd1417,16'd1944,-16'd6209,-16'd5192,-16'd8364,-16'd1295,-16'd4058,16'd73};
dout[954]={ -16'd6910,16'd6087,-16'd3347,-16'd1886,-16'd5504,16'd211,16'd8933,16'd7066,16'd6229,-16'd5779,-16'd4359,-16'd1691,-16'd1004,16'd6116,-16'd4357,16'd4921,-16'd7644,16'd6135,16'd5989,-16'd7033,16'd5756,16'd2952,-16'd2586,-16'd1470,-16'd604,16'd5930,16'd4780,-16'd4457,16'd6091,16'd508,-16'd3450,16'd6093,16'd3096,16'd4655,-16'd8611,-16'd779};
dout[955]={ -16'd5002,16'd6343,-16'd4708,-16'd3749,16'd5006,16'd1156,16'd2486,16'd1614,-16'd3578,-16'd8011,16'd1368,-16'd5311,-16'd697,16'd2219,-16'd3138,16'd427,-16'd4596,16'd5159,16'd4195,-16'd1593,-16'd1044,-16'd6643,-16'd2775,-16'd1414,-16'd1870,16'd1653,-16'd2577,16'd1657,16'd4267,16'd4653,-16'd3950,-16'd3263,16'd5451,-16'd124,-16'd2608,-16'd9287};
dout[956]={ -16'd7229,16'd6320,-16'd8310,16'd2669,16'd5150,-16'd3733,16'd6428,16'd466,-16'd6473,-16'd417,16'd6085,16'd2611,-16'd6915,16'd6613,-16'd2532,-16'd7150,-16'd4677,16'd3776,-16'd6650,-16'd7009,-16'd1014,-16'd3826,-16'd4299,16'd4259,-16'd2785,16'd1631,-16'd3006,-16'd5852,16'd3038,-16'd3756,16'd7958,-16'd733,-16'd4829,-16'd3386,-16'd5428,16'd317};
dout[957]={ -16'd8581,-16'd3444,-16'd4001,16'd1128,16'd3656,-16'd7281,-16'd2310,16'd2799,16'd1812,-16'd1521,16'd7179,-16'd2882,-16'd7190,16'd5740,-16'd6957,-16'd6783,-16'd8549,16'd4790,-16'd4631,16'd2994,-16'd1637,-16'd3892,16'd4659,-16'd6878,16'd6267,-16'd5052,-16'd5062,16'd5891,16'd2011,-16'd6333,16'd1187,-16'd3756,-16'd5031,16'd985,16'd6573,16'd5580};
dout[958]={ -16'd4137,16'd6254,-16'd203,16'd3721,16'd4754,-16'd7393,-16'd1234,16'd6334,16'd2019,-16'd6098,-16'd2467,16'd4641,16'd1795,-16'd403,16'd3823,16'd5671,-16'd1605,16'd7351,-16'd7924,16'd2494,16'd3560,16'd5127,-16'd1609,16'd1621,-16'd1135,16'd663,16'd813,16'd5920,16'd6334,-16'd3955,-16'd2603,-16'd5240,-16'd7068,-16'd2175,-16'd6973,-16'd2833};
dout[959]={ 16'd3649,-16'd5170,16'd4859,16'd4115,16'd3170,-16'd4270,-16'd5784,-16'd2761,-16'd2848,-16'd5127,16'd3078,-16'd87,16'd5546,16'd4977,16'd1917,16'd1312,16'd1060,16'd160,-16'd2609,16'd1643,16'd2815,-16'd1036,-16'd341,16'd3014,16'd7997,-16'd8315,16'd41,16'd5676,-16'd6855,16'd2402,-16'd5772,16'd6996,16'd6257,-16'd1780,16'd5037,-16'd3822};
dout[960]={ -16'd1824,16'd13690,-16'd5062,-16'd5217,-16'd929,16'd7376,16'd3790,16'd2020,-16'd8245,16'd463,-16'd4681,-16'd1142,-16'd1833,-16'd140,-16'd1108,16'd1370,16'd2087,16'd93,-16'd10207,16'd1349,-16'd2918,16'd5001,-16'd1953,16'd3063,16'd6443,-16'd4995,16'd317,-16'd8647,16'd3883,-16'd3284,16'd2755,16'd6070,16'd3696,-16'd10369,-16'd236,16'd1044};
dout[961]={ -16'd2851,16'd7250,16'd1905,-16'd954,-16'd5652,16'd4734,16'd2627,16'd5243,-16'd6844,16'd3740,16'd3274,16'd9206,16'd3179,-16'd5032,16'd3501,16'd1141,16'd4674,-16'd1113,16'd49,16'd4126,-16'd3415,-16'd30,-16'd3383,16'd6529,16'd6159,-16'd6324,16'd3067,-16'd5967,16'd5981,16'd7581,16'd727,16'd1070,-16'd4059,16'd413,-16'd8929,-16'd1307};
dout[962]={ 16'd1125,16'd4062,16'd7178,-16'd3518,-16'd8460,-16'd1179,16'd2713,-16'd8105,-16'd3419,16'd3819,-16'd7920,16'd834,16'd3562,16'd9739,-16'd7313,16'd3694,-16'd7233,16'd2884,-16'd6575,16'd2936,16'd6138,-16'd859,16'd1553,16'd1234,16'd2631,-16'd2474,-16'd1252,-16'd979,-16'd6519,-16'd642,-16'd3198,-16'd3130,16'd1945,-16'd445,16'd1163,-16'd8836};
dout[963]={ -16'd703,16'd1178,16'd8504,-16'd9085,16'd2299,16'd6040,16'd6413,16'd6324,-16'd2308,-16'd3025,-16'd7145,16'd3184,-16'd7567,-16'd1052,16'd5359,-16'd6825,16'd6184,-16'd1087,16'd3893,-16'd11402,16'd1253,16'd274,16'd2369,16'd6922,-16'd6459,16'd3159,-16'd80,-16'd4119,16'd1144,-16'd2379,-16'd9770,16'd4634,-16'd4333,-16'd4914,-16'd4133,-16'd6203};
dout[964]={ -16'd1433,-16'd2605,-16'd1170,16'd2511,16'd1412,-16'd3589,16'd2153,-16'd1421,16'd6908,16'd5655,16'd5066,16'd816,16'd7523,-16'd9884,16'd4857,-16'd2842,16'd93,16'd6047,16'd6674,-16'd8164,16'd1183,16'd6466,16'd5443,16'd3479,-16'd3547,-16'd2093,-16'd3562,16'd1232,16'd876,-16'd1912,16'd2544,-16'd6655,16'd2490,16'd2028,-16'd410,-16'd3387};
dout[965]={ 16'd5437,16'd7887,16'd623,-16'd4775,-16'd3200,16'd1681,16'd3133,16'd3278,-16'd2103,-16'd7639,16'd3456,-16'd6155,16'd4148,-16'd2258,16'd1243,-16'd5810,16'd786,-16'd10,-16'd10236,-16'd2191,-16'd6739,16'd5766,16'd4017,-16'd4544,-16'd77,16'd225,-16'd789,16'd340,16'd4407,16'd3741,-16'd1246,16'd6247,-16'd7424,16'd2633,16'd4950,-16'd9112};
dout[966]={ 16'd1293,-16'd1013,-16'd2313,-16'd7373,-16'd5430,-16'd4582,-16'd3581,-16'd665,-16'd2093,-16'd5052,-16'd3153,-16'd3487,16'd2901,-16'd1780,-16'd3599,-16'd61,-16'd7636,-16'd585,-16'd5502,16'd1961,16'd2984,16'd915,16'd5693,-16'd356,16'd8242,16'd5135,16'd5461,16'd1803,-16'd2117,-16'd3193,16'd103,-16'd3301,-16'd7151,16'd5413,16'd2518,16'd7360};
dout[967]={ -16'd2319,16'd2450,16'd3370,16'd4256,-16'd1311,16'd2219,16'd3208,-16'd3876,-16'd992,16'd597,16'd2048,16'd5002,16'd468,16'd5932,16'd4623,-16'd2535,-16'd2895,16'd3179,-16'd2861,-16'd568,-16'd5885,-16'd3817,-16'd3869,16'd4152,16'd5569,-16'd4977,16'd4738,16'd9289,-16'd1438,16'd3558,-16'd5776,-16'd6263,-16'd8357,-16'd4634,-16'd1863,-16'd3114};
dout[968]={ 16'd4665,16'd183,16'd360,-16'd7755,-16'd2222,16'd4376,16'd3701,16'd8947,-16'd579,-16'd2009,16'd3091,16'd118,16'd1824,16'd5453,16'd4243,-16'd3867,16'd5730,16'd2002,-16'd3680,16'd4773,16'd2184,-16'd1834,-16'd2374,16'd3163,-16'd4760,-16'd2063,16'd2182,-16'd2154,-16'd806,-16'd5410,-16'd5527,-16'd4545,16'd3743,16'd8016,-16'd1675,16'd8713};
dout[969]={ -16'd6991,16'd6409,16'd6284,-16'd5271,16'd4328,-16'd4740,16'd4558,16'd616,16'd6931,-16'd1544,16'd2569,-16'd3538,-16'd5461,16'd3370,-16'd7764,-16'd1328,-16'd4107,16'd5349,-16'd5348,-16'd4635,16'd2885,16'd5534,-16'd4286,-16'd2850,-16'd5468,-16'd10221,-16'd6358,16'd7655,-16'd1825,-16'd4458,16'd5683,-16'd6795,-16'd6960,-16'd2826,-16'd2008,16'd9016};
dout[970]={ 16'd2983,16'd1658,16'd4986,16'd5741,16'd907,16'd2827,16'd8801,-16'd6367,-16'd1439,-16'd3631,16'd5781,16'd2869,-16'd3836,16'd7844,16'd845,-16'd6020,16'd1251,16'd7390,-16'd2398,16'd3054,16'd3861,16'd2594,16'd3228,16'd1614,-16'd13171,-16'd5349,16'd4016,-16'd996,-16'd2242,16'd4598,16'd6287,-16'd5486,16'd1285,-16'd12395,-16'd1906,-16'd13522};
dout[971]={ 16'd9568,-16'd2794,-16'd413,16'd6470,16'd831,-16'd4942,16'd1366,16'd95,16'd2449,-16'd2734,16'd3781,16'd3446,16'd2925,16'd6976,-16'd2938,-16'd8062,-16'd9660,-16'd1614,16'd3209,16'd5198,16'd4927,-16'd1141,-16'd6163,-16'd2728,16'd217,-16'd8851,-16'd758,-16'd8755,16'd1612,16'd484,-16'd1322,16'd5995,16'd2688,-16'd5306,-16'd1401,16'd3006};
dout[972]={ -16'd3286,-16'd791,-16'd244,-16'd1973,-16'd4023,-16'd7997,16'd3474,-16'd7113,-16'd485,16'd2566,-16'd6361,-16'd3246,-16'd11745,16'd6612,-16'd9390,-16'd3824,-16'd2457,-16'd2382,16'd3352,16'd836,-16'd373,-16'd5181,16'd8127,-16'd4876,16'd8552,16'd4522,-16'd1013,-16'd3777,16'd1160,16'd7235,16'd2542,-16'd4520,-16'd8051,-16'd4100,16'd651,-16'd11219};
dout[973]={ -16'd5158,16'd1154,16'd5579,-16'd422,-16'd4359,16'd3089,-16'd6696,16'd2319,16'd5289,16'd417,-16'd1421,-16'd7252,16'd1631,-16'd3287,-16'd4350,-16'd397,16'd5483,-16'd3681,-16'd2544,-16'd5505,-16'd6601,-16'd5231,16'd4594,16'd4537,-16'd7772,-16'd2765,-16'd5398,16'd2094,16'd3554,16'd3373,-16'd12221,-16'd2661,-16'd8833,16'd5064,16'd6198,-16'd3144};
dout[974]={ 16'd4968,16'd8863,-16'd5121,-16'd4873,-16'd2588,-16'd2379,-16'd3820,-16'd1959,16'd7577,16'd5487,-16'd3261,-16'd460,-16'd7132,-16'd700,-16'd243,-16'd1805,-16'd730,16'd63,-16'd3929,-16'd4426,16'd6811,16'd3483,-16'd8781,16'd1464,-16'd4719,16'd6054,-16'd7348,16'd6752,16'd7734,16'd1074,16'd792,16'd6376,-16'd4815,-16'd958,-16'd6375,-16'd8613};
dout[975]={ -16'd2741,16'd5967,16'd3455,-16'd3990,16'd3624,16'd3294,16'd1248,-16'd26,-16'd84,-16'd926,-16'd1384,-16'd6537,16'd5662,-16'd1382,16'd3839,-16'd4793,16'd6834,-16'd2123,-16'd7286,-16'd834,16'd5369,16'd458,-16'd5911,16'd2666,16'd4007,-16'd4006,-16'd8070,-16'd272,16'd3896,-16'd5880,16'd4305,16'd6300,16'd3216,-16'd1719,-16'd75,-16'd2648};
dout[976]={ 16'd1697,-16'd5222,16'd2379,-16'd7709,-16'd8006,16'd7540,16'd6902,-16'd2415,-16'd59,16'd3218,16'd2128,16'd5627,-16'd8785,-16'd3335,16'd2797,16'd5311,-16'd1354,16'd3159,-16'd4817,-16'd3691,16'd2811,-16'd2276,-16'd5552,16'd1722,-16'd3944,16'd1057,16'd2797,16'd539,16'd2833,16'd3684,-16'd3400,-16'd547,16'd4199,-16'd8311,-16'd4861,-16'd2924};
dout[977]={ 16'd3584,16'd1933,16'd1002,-16'd2269,16'd6156,16'd3561,16'd3882,16'd7966,16'd5901,-16'd108,16'd2341,-16'd5896,-16'd228,16'd6142,16'd1403,16'd1072,16'd4676,16'd1379,-16'd3348,16'd6484,16'd5802,-16'd5756,16'd4167,-16'd3299,-16'd4432,-16'd5120,-16'd732,16'd2471,16'd432,16'd3538,16'd2793,-16'd736,-16'd7979,-16'd4036,-16'd3114,-16'd4380};
dout[978]={ 16'd2280,16'd5510,16'd4881,-16'd951,-16'd2632,16'd5783,16'd4958,16'd6754,-16'd6531,-16'd5252,16'd7206,-16'd6024,16'd237,16'd2145,-16'd7944,-16'd2254,16'd1233,-16'd1236,16'd268,16'd4117,16'd330,-16'd6548,16'd3503,-16'd4026,-16'd268,16'd2602,-16'd7450,16'd9026,16'd6307,16'd703,16'd698,-16'd84,16'd67,16'd4001,-16'd5668,-16'd3814};
dout[979]={ -16'd2322,-16'd2824,-16'd1952,16'd4546,-16'd7405,-16'd3951,-16'd4544,-16'd4922,16'd699,-16'd6113,16'd2066,-16'd4591,-16'd3159,16'd2787,-16'd6360,16'd1304,-16'd2794,16'd4408,16'd7293,-16'd5691,16'd737,-16'd2120,16'd1814,-16'd2587,16'd7232,16'd2495,-16'd8113,16'd146,-16'd6755,-16'd1808,-16'd4758,-16'd3484,-16'd7271,16'd4113,16'd2899,16'd3451};
dout[980]={ 16'd2892,16'd3206,16'd6520,16'd1814,-16'd165,16'd3598,16'd5724,-16'd5728,-16'd1675,16'd2966,-16'd2859,-16'd235,16'd4751,16'd494,-16'd9264,-16'd7125,16'd305,16'd9271,-16'd4063,-16'd327,16'd8,-16'd4748,16'd106,-16'd74,-16'd9127,-16'd1405,16'd6836,-16'd6773,-16'd7707,16'd3040,-16'd1868,-16'd717,16'd4306,-16'd12465,16'd382,16'd5607};
dout[981]={ 16'd5337,-16'd9629,-16'd1312,-16'd4175,-16'd354,16'd6095,16'd8224,16'd716,-16'd4576,16'd5021,16'd1190,16'd11155,-16'd7099,-16'd1725,16'd1421,16'd4454,16'd5398,16'd1165,16'd6345,16'd6389,16'd4534,16'd820,16'd7020,16'd6737,16'd1790,16'd2680,16'd955,-16'd8339,-16'd2257,-16'd1765,16'd2629,-16'd5148,-16'd1368,-16'd7447,-16'd4593,16'd2455};
dout[982]={ 16'd876,-16'd8593,16'd1992,-16'd5775,16'd440,16'd914,16'd383,-16'd12388,-16'd204,-16'd1196,-16'd1053,16'd4124,-16'd5579,16'd4994,16'd1296,16'd2440,16'd1784,-16'd3412,16'd6871,16'd9124,16'd7301,16'd5275,-16'd948,-16'd2820,-16'd1576,16'd349,16'd10709,16'd506,16'd4688,-16'd1912,16'd2125,-16'd2485,-16'd9459,-16'd1322,16'd3237,-16'd11936};
dout[983]={ 16'd5975,-16'd1139,16'd2026,-16'd313,-16'd2139,-16'd618,-16'd6224,-16'd2774,-16'd5949,16'd573,16'd2053,16'd1739,-16'd8297,16'd1392,-16'd3827,16'd825,-16'd3502,16'd2743,16'd1914,-16'd10147,16'd1822,16'd328,16'd1024,16'd1729,16'd5469,16'd4794,-16'd7856,-16'd1457,16'd1417,-16'd1640,-16'd5928,-16'd2206,-16'd4504,-16'd2391,-16'd2526,-16'd5570};
dout[984]={ 16'd1626,-16'd6900,16'd4880,-16'd10542,-16'd1604,16'd6393,-16'd6741,16'd6772,-16'd3923,-16'd1654,16'd3346,-16'd5881,-16'd10378,-16'd14756,-16'd6618,16'd2190,16'd6084,16'd6383,-16'd609,-16'd2319,16'd2616,-16'd2568,16'd1514,16'd1836,-16'd9616,-16'd5678,-16'd2453,16'd6332,-16'd3853,-16'd925,-16'd8751,-16'd4818,16'd2524,16'd5111,16'd6341,-16'd8805};
dout[985]={ -16'd1292,-16'd6671,-16'd987,-16'd1825,16'd4598,16'd2345,-16'd2484,16'd4710,16'd1653,16'd2165,16'd1736,-16'd186,16'd1309,-16'd6076,16'd3629,16'd379,16'd6092,-16'd7622,-16'd2071,16'd775,16'd3793,-16'd262,16'd5907,-16'd5054,-16'd8429,16'd2072,16'd1588,16'd3965,-16'd1031,16'd5557,-16'd1368,-16'd4058,-16'd1879,16'd4298,16'd938,-16'd242};
dout[986]={ 16'd932,16'd439,-16'd8429,16'd183,16'd1359,16'd1666,16'd4456,-16'd2676,16'd6137,-16'd3726,-16'd4738,-16'd5005,-16'd1668,16'd1010,-16'd3959,16'd1428,16'd5598,16'd1274,-16'd6559,-16'd2023,16'd4094,-16'd101,-16'd4512,-16'd2166,-16'd824,-16'd5349,-16'd3221,-16'd3974,-16'd6731,-16'd1564,-16'd1310,-16'd2371,16'd3492,16'd1878,16'd1280,-16'd4214};
dout[987]={ 16'd4684,-16'd5903,16'd1953,-16'd4017,16'd423,16'd1940,-16'd4124,16'd3524,-16'd3209,16'd1948,16'd2222,-16'd482,-16'd2678,-16'd5852,-16'd4941,16'd2289,-16'd3315,16'd5879,-16'd2939,16'd3025,-16'd8312,16'd6722,-16'd3153,-16'd7552,16'd3889,16'd2630,16'd7907,16'd542,16'd4078,-16'd4494,-16'd4156,16'd3655,-16'd6921,-16'd241,-16'd6111,16'd3116};
dout[988]={ -16'd1918,16'd1296,16'd44,-16'd5312,-16'd2534,16'd2150,16'd484,-16'd5582,16'd967,16'd713,16'd6204,16'd4323,-16'd6189,-16'd6783,16'd2180,-16'd6807,-16'd5788,16'd824,16'd187,-16'd5055,-16'd283,16'd1321,16'd1574,-16'd1183,16'd2010,-16'd8131,-16'd1715,16'd1526,-16'd3739,16'd2310,16'd3423,-16'd7231,-16'd644,-16'd2764,-16'd3872,16'd1357};
dout[989]={ 16'd1877,16'd2566,16'd4799,-16'd2321,16'd4562,16'd2566,-16'd6793,-16'd4455,16'd5277,16'd2708,16'd6576,-16'd958,16'd181,-16'd5427,-16'd8549,16'd4493,-16'd2368,16'd4594,16'd10855,16'd5966,16'd5556,-16'd5105,16'd7135,-16'd7816,16'd3837,16'd3751,-16'd1662,16'd8059,16'd2251,16'd281,-16'd8010,-16'd1731,-16'd2738,16'd151,16'd8344,16'd6639};
dout[990]={ -16'd862,-16'd68,-16'd1011,-16'd662,-16'd5286,-16'd3919,16'd2787,-16'd1937,-16'd10842,-16'd1441,-16'd158,16'd1076,-16'd3408,16'd11832,-16'd6978,-16'd4061,16'd3305,16'd8215,16'd5657,16'd1517,-16'd500,-16'd8878,16'd5883,16'd6057,-16'd6000,16'd7409,16'd330,16'd3070,16'd4571,-16'd891,16'd3950,16'd6815,16'd3017,-16'd829,16'd8234,16'd1929};
dout[991]={ -16'd7436,-16'd557,-16'd4426,-16'd1849,-16'd3897,-16'd6872,16'd2080,-16'd12924,-16'd633,16'd265,16'd6715,16'd5867,-16'd11787,16'd8675,16'd1275,-16'd3705,16'd7125,16'd835,16'd6232,-16'd44,-16'd4811,16'd4429,-16'd511,16'd8343,-16'd1463,-16'd2340,-16'd1153,-16'd4107,16'd712,16'd4768,16'd6624,-16'd5266,-16'd7917,16'd4856,16'd1845,-16'd3270};
dout[992]={ 16'd3960,-16'd3163,16'd7030,-16'd1654,16'd2353,16'd3944,-16'd2113,-16'd5801,-16'd12242,16'd5298,-16'd4954,16'd4824,-16'd5467,16'd5987,-16'd3063,-16'd2530,16'd5297,16'd7116,16'd6174,-16'd3445,-16'd2344,-16'd6066,16'd4144,16'd10010,-16'd4108,16'd2328,-16'd3016,-16'd4780,-16'd2401,16'd1655,16'd6566,16'd3960,-16'd8989,16'd5045,16'd6414,-16'd6319};
dout[993]={ -16'd3993,16'd3170,-16'd3619,-16'd393,16'd3361,-16'd3253,-16'd13757,-16'd8190,-16'd1215,16'd2548,-16'd8674,-16'd1683,-16'd3703,-16'd8206,16'd4299,-16'd6001,16'd6461,-16'd2497,16'd3515,-16'd3196,16'd5562,-16'd5887,-16'd4694,16'd1727,16'd4624,-16'd663,-16'd8628,-16'd526,-16'd1626,16'd2024,-16'd11128,-16'd2337,-16'd6220,16'd847,-16'd1637,16'd6615};
dout[994]={ -16'd1898,-16'd5569,16'd7008,-16'd6117,-16'd1305,-16'd2341,-16'd1379,-16'd5190,-16'd6986,-16'd5336,-16'd2193,-16'd5940,16'd4355,-16'd5692,16'd4317,-16'd4316,-16'd4008,16'd2532,16'd4146,16'd2823,-16'd4440,-16'd1391,-16'd2653,16'd8490,-16'd3688,-16'd394,-16'd9129,-16'd2097,-16'd1096,-16'd2154,16'd3871,-16'd9766,-16'd2752,16'd1584,-16'd5318,16'd4551};
dout[995]={ -16'd1374,-16'd5469,-16'd5025,-16'd3215,16'd264,-16'd2590,16'd6024,-16'd853,16'd7651,16'd8442,-16'd8578,-16'd4904,-16'd7694,-16'd5039,-16'd8684,-16'd2991,16'd834,-16'd3822,-16'd6171,-16'd1843,-16'd4092,16'd705,16'd4792,-16'd1416,16'd1308,-16'd3944,16'd471,-16'd3780,16'd3102,-16'd1165,16'd2560,-16'd1476,16'd6,-16'd2920,-16'd2538,-16'd1501};
dout[996]={ 16'd1490,-16'd7164,16'd2958,-16'd10360,16'd5773,-16'd6846,-16'd6429,16'd5028,16'd1412,-16'd2135,16'd5753,-16'd4129,-16'd7675,16'd7200,16'd4308,-16'd8021,-16'd773,-16'd4187,16'd4964,-16'd2145,-16'd414,16'd2701,-16'd4052,-16'd4557,16'd2225,16'd7738,16'd4316,-16'd3296,16'd907,16'd1637,16'd3089,16'd2740,16'd2828,16'd2642,-16'd2643,16'd4372};
dout[997]={ -16'd4053,-16'd1184,-16'd1329,-16'd9452,16'd2618,16'd1753,16'd4334,16'd4949,16'd5030,-16'd2530,16'd5139,-16'd5752,-16'd2882,-16'd1964,16'd2544,16'd5691,16'd2415,16'd1760,16'd2978,16'd4124,-16'd2396,16'd3791,16'd3167,-16'd6182,16'd4042,16'd527,16'd748,-16'd2989,16'd1232,16'd4059,-16'd4898,-16'd5474,-16'd4495,16'd3076,-16'd3666,16'd4126};
dout[998]={ -16'd5673,16'd3068,-16'd1296,16'd2889,-16'd3878,16'd4554,-16'd422,-16'd2141,16'd3200,-16'd5621,-16'd3081,-16'd7225,-16'd135,-16'd6177,-16'd9892,-16'd9236,16'd3048,-16'd467,-16'd3330,16'd666,16'd146,16'd2539,-16'd5793,16'd4100,16'd4311,-16'd7104,-16'd2485,16'd5671,16'd4227,-16'd1697,16'd2507,16'd2569,16'd525,16'd5485,-16'd1834,16'd87};
dout[999]={ -16'd1957,-16'd3190,-16'd4637,16'd2157,16'd2310,-16'd3473,-16'd3253,-16'd2811,-16'd2429,-16'd1551,-16'd4918,-16'd3149,-16'd5496,16'd1845,16'd845,-16'd6464,-16'd2280,-16'd3372,16'd2996,-16'd910,-16'd3140,-16'd3315,-16'd3861,-16'd2712,-16'd207,-16'd8061,-16'd8003,16'd6167,16'd3290,-16'd3351,-16'd911,16'd511,16'd5103,16'd5709,-16'd4576,16'd5941};
dout[1000]={ 16'd53,-16'd15600,16'd0,16'd7287,-16'd1429,16'd6335,16'd5135,-16'd3053,-16'd10224,16'd1032,-16'd8708,16'd404,-16'd4272,16'd6642,-16'd1930,-16'd9052,-16'd6921,16'd2165,-16'd1637,16'd1743,-16'd4338,16'd1901,16'd2534,-16'd5958,-16'd12261,16'd5683,16'd4594,16'd2970,-16'd4921,16'd1557,16'd5941,-16'd1675,16'd1482,-16'd8435,16'd8912,16'd9179};
dout[1001]={ -16'd3444,-16'd7352,16'd1876,-16'd3040,-16'd1430,16'd1750,16'd7735,16'd4750,-16'd8806,16'd4353,-16'd7860,16'd3148,-16'd2234,16'd6561,-16'd3999,-16'd456,-16'd8501,-16'd402,16'd2437,-16'd866,16'd3467,-16'd2510,16'd5172,16'd7808,-16'd1737,-16'd735,16'd736,-16'd9358,-16'd6534,-16'd2815,16'd4208,16'd2589,16'd1527,16'd753,-16'd2935,16'd8128};
dout[1002]={ 16'd317,-16'd2787,16'd6080,16'd41,16'd1018,-16'd8745,-16'd8600,16'd6952,-16'd6496,-16'd8047,-16'd9453,16'd10329,16'd3604,16'd10457,-16'd7389,-16'd3258,16'd2506,16'd5029,16'd3252,-16'd195,-16'd4097,16'd3547,16'd6428,-16'd4371,16'd2909,16'd7933,16'd7491,-16'd5887,-16'd1048,-16'd1772,-16'd5181,-16'd8479,16'd4350,16'd6610,-16'd1103,-16'd3315};
dout[1003]={ -16'd3840,-16'd7086,-16'd4959,16'd1986,-16'd4108,16'd3517,-16'd3791,-16'd5762,-16'd5642,16'd3363,-16'd6056,-16'd2720,16'd3725,-16'd9934,16'd2628,-16'd6189,16'd3001,-16'd3122,16'd3481,-16'd13479,-16'd9310,-16'd3349,16'd850,16'd7121,16'd1617,16'd1525,-16'd12044,16'd208,-16'd8409,16'd2433,-16'd13310,16'd2200,16'd336,16'd2767,-16'd7112,16'd2808};
dout[1004]={ -16'd756,16'd1027,-16'd6474,-16'd8330,-16'd364,-16'd1350,-16'd5774,-16'd6436,16'd409,-16'd1788,16'd4424,-16'd4087,16'd6000,-16'd5834,-16'd5862,-16'd4099,-16'd5369,-16'd2732,16'd5032,16'd1410,-16'd3123,-16'd4479,-16'd5888,16'd3901,16'd2419,16'd5073,-16'd11076,16'd9268,-16'd282,-16'd2965,-16'd7962,16'd330,-16'd312,16'd1930,16'd873,-16'd3188};
dout[1005]={ 16'd5568,-16'd4772,16'd4905,-16'd6254,-16'd1015,16'd5313,-16'd3068,16'd5351,-16'd1277,16'd9338,-16'd4016,-16'd6423,16'd4416,-16'd4019,16'd788,-16'd1269,16'd3416,-16'd951,16'd1531,16'd1960,-16'd6188,-16'd3697,-16'd8486,-16'd363,16'd403,16'd2772,16'd353,-16'd3209,16'd5158,-16'd833,-16'd6843,-16'd880,-16'd9245,16'd7394,16'd798,16'd4279};
dout[1006]={ -16'd5538,16'd3086,16'd1828,-16'd11408,16'd3936,-16'd1212,-16'd3630,-16'd6593,-16'd1824,16'd7574,16'd5903,16'd548,-16'd1083,-16'd3976,-16'd2565,-16'd802,16'd3422,16'd4914,16'd1166,-16'd2266,-16'd6245,-16'd6905,-16'd2235,-16'd5760,16'd4952,16'd1090,-16'd2074,16'd4488,16'd2154,-16'd1632,16'd4405,16'd5554,16'd1671,-16'd147,16'd1807,-16'd5831};
dout[1007]={ -16'd3424,16'd2520,16'd3916,-16'd4542,16'd143,-16'd6789,-16'd1026,-16'd1739,16'd2705,16'd4826,16'd4369,-16'd2765,-16'd2451,-16'd3434,16'd4198,16'd4751,16'd372,-16'd4730,16'd4945,16'd4912,16'd3020,16'd2315,-16'd3650,-16'd4541,-16'd943,-16'd3016,-16'd398,-16'd4392,-16'd5058,-16'd4400,-16'd8980,-16'd9677,16'd5494,16'd2030,-16'd7937,16'd2546};
dout[1008]={ -16'd6748,16'd6075,16'd5545,-16'd10772,16'd5532,16'd3668,-16'd4735,16'd6002,16'd6872,16'd5179,-16'd4587,-16'd2844,-16'd5251,-16'd1451,16'd3466,-16'd6314,-16'd8987,16'd5356,16'd691,-16'd5462,16'd425,16'd2745,16'd6062,-16'd3646,16'd6543,16'd6617,16'd2451,16'd1985,16'd7720,-16'd7988,16'd868,16'd2933,16'd2283,-16'd2184,-16'd6357,16'd4867};
dout[1009]={ -16'd1568,-16'd3947,-16'd6073,-16'd4805,16'd4724,-16'd6977,-16'd1554,-16'd6627,-16'd164,-16'd8634,16'd79,16'd3250,-16'd4388,16'd4484,-16'd3927,-16'd6812,16'd6156,16'd7177,16'd2391,16'd4559,-16'd1096,16'd316,16'd7236,16'd3020,16'd3859,-16'd3612,16'd2826,16'd4638,-16'd2425,-16'd8159,-16'd5573,-16'd1040,-16'd2766,-16'd2643,16'd51,-16'd4832};
dout[1010]={ -16'd8257,-16'd2255,16'd179,16'd6252,16'd1840,16'd6289,-16'd4668,-16'd103,-16'd3687,-16'd3432,-16'd7558,16'd6463,-16'd1063,-16'd1475,-16'd3862,16'd5597,16'd3506,-16'd6879,16'd7286,16'd7109,-16'd2713,-16'd719,-16'd3751,16'd4486,16'd3847,16'd13263,16'd9223,16'd9005,-16'd4019,-16'd4673,16'd5140,-16'd4089,16'd3092,-16'd2006,-16'd5667,16'd7667};
dout[1011]={ -16'd10411,16'd1308,-16'd2583,-16'd1006,16'd4500,16'd73,-16'd3909,-16'd6669,16'd7103,-16'd5563,-16'd7691,16'd12326,16'd267,16'd4532,-16'd5546,16'd3917,16'd465,16'd8415,-16'd2941,16'd4831,16'd465,16'd3799,-16'd7936,16'd1050,16'd2337,16'd9709,-16'd287,16'd3553,-16'd1122,16'd2049,16'd5214,-16'd2811,16'd3906,16'd8250,16'd3835,-16'd2069};
dout[1012]={ -16'd6342,-16'd2786,16'd4907,-16'd2041,16'd490,-16'd7276,-16'd4987,16'd5180,-16'd8734,-16'd1967,-16'd5184,16'd6596,-16'd7085,16'd3371,-16'd3387,-16'd1736,16'd2518,16'd2535,-16'd2598,16'd1037,-16'd1725,-16'd2737,-16'd4112,16'd5868,16'd3682,16'd5262,16'd1620,-16'd5883,-16'd2323,-16'd4323,16'd2641,-16'd7187,16'd2050,-16'd3805,16'd651,16'd5678};
dout[1013]={ -16'd1229,-16'd3675,16'd550,-16'd754,-16'd6652,16'd4823,-16'd10524,16'd617,-16'd5550,16'd4185,-16'd110,-16'd2087,16'd2354,-16'd5803,-16'd8159,-16'd6369,16'd224,-16'd142,16'd8215,-16'd902,-16'd8568,16'd1356,-16'd5821,-16'd4630,-16'd4091,16'd1805,-16'd12370,-16'd958,16'd4454,-16'd4581,-16'd13485,16'd145,-16'd7869,16'd774,-16'd1982,16'd1602};
dout[1014]={ -16'd5842,-16'd1330,16'd4800,16'd1499,-16'd4428,16'd2726,-16'd11923,-16'd22,-16'd4470,16'd7110,16'd5040,-16'd3403,16'd7205,16'd1807,-16'd5117,16'd4523,16'd250,-16'd997,-16'd6210,16'd95,-16'd7819,16'd681,16'd519,16'd4834,-16'd2893,16'd737,-16'd8849,16'd5768,-16'd1746,-16'd8008,-16'd4190,-16'd7568,16'd1462,16'd3459,-16'd6737,-16'd6401};
dout[1015]={ 16'd6489,-16'd885,16'd5970,-16'd10375,-16'd7763,-16'd5648,16'd1752,-16'd4185,-16'd2691,-16'd2053,16'd3121,-16'd2798,16'd1437,-16'd3546,-16'd6619,-16'd6522,-16'd3177,-16'd3134,16'd7772,16'd7300,-16'd1296,-16'd7602,16'd2497,-16'd2608,-16'd1555,16'd3859,-16'd8614,16'd3944,-16'd6752,-16'd2801,-16'd405,-16'd756,-16'd1058,-16'd3761,16'd3794,16'd5166};
dout[1016]={ -16'd473,-16'd4181,16'd327,-16'd10270,16'd2674,16'd2880,-16'd8239,-16'd9210,16'd394,-16'd1359,-16'd7211,16'd2444,-16'd3936,-16'd6010,-16'd1827,-16'd1555,-16'd8022,16'd1641,-16'd6176,-16'd5715,-16'd74,16'd1611,16'd5607,16'd792,-16'd112,-16'd1514,-16'd708,-16'd2479,16'd953,-16'd4822,16'd4432,-16'd1263,-16'd4282,-16'd1584,-16'd2821,16'd3019};
dout[1017]={ -16'd1921,-16'd3992,16'd1588,-16'd8039,16'd1055,16'd4582,16'd6708,16'd5794,-16'd582,-16'd1100,-16'd139,16'd49,-16'd5307,-16'd3554,16'd316,-16'd193,-16'd7515,-16'd3774,16'd3696,16'd5702,-16'd5531,-16'd4588,-16'd5619,-16'd3284,16'd6469,16'd1610,16'd7219,16'd4302,16'd4034,-16'd2997,16'd4131,16'd3111,16'd2455,16'd17,-16'd2824,16'd5173};
dout[1018]={ -16'd6442,16'd4431,16'd416,-16'd6299,-16'd4953,-16'd4669,16'd924,-16'd4898,-16'd2844,-16'd2214,16'd3952,-16'd6657,-16'd3576,-16'd5311,16'd4876,-16'd39,-16'd255,-16'd3976,16'd3287,-16'd5226,-16'd1511,-16'd7398,-16'd2929,16'd4127,-16'd3048,-16'd1253,16'd5667,-16'd3232,16'd7844,-16'd572,16'd5432,-16'd9649,16'd5581,16'd4727,16'd5616,16'd481};
dout[1019]={ -16'd1019,-16'd2354,16'd2585,-16'd9564,16'd1845,-16'd9572,16'd1363,-16'd8632,16'd6760,16'd4192,16'd5506,-16'd4381,16'd4309,16'd1526,16'd4850,16'd72,-16'd6721,-16'd1238,-16'd3165,-16'd2614,16'd7324,16'd2964,-16'd2193,-16'd3970,16'd1398,-16'd2648,-16'd7648,-16'd4566,-16'd466,-16'd1259,16'd182,16'd1045,-16'd5922,-16'd2326,-16'd2495,-16'd4245};
dout[1020]={ -16'd4715,-16'd4535,-16'd8843,16'd482,-16'd2962,-16'd2905,-16'd7913,16'd2915,-16'd3839,-16'd476,16'd2328,-16'd2842,-16'd4664,16'd858,-16'd1089,16'd8657,-16'd5656,16'd4253,16'd6984,16'd8748,-16'd91,16'd4251,-16'd518,16'd4170,-16'd871,16'd7922,16'd3147,16'd1983,16'd2861,-16'd4740,-16'd5141,16'd1965,16'd5906,16'd1129,-16'd3331,-16'd2622};
dout[1021]={ -16'd4473,-16'd2144,-16'd1637,16'd3267,16'd2124,16'd6564,-16'd2938,-16'd2263,16'd5699,-16'd8395,-16'd3838,16'd4968,-16'd569,16'd2224,-16'd473,-16'd2978,16'd2460,-16'd4524,-16'd2789,16'd7549,-16'd6036,-16'd8291,-16'd5630,-16'd7450,16'd5319,16'd10066,16'd5856,16'd5527,-16'd6558,16'd4772,16'd3889,-16'd5031,-16'd2080,-16'd2870,-16'd6807,16'd2567};
dout[1022]={ 16'd1934,-16'd6307,16'd8942,16'd6028,16'd408,16'd4157,-16'd8930,16'd6925,-16'd6619,-16'd3966,16'd3298,-16'd1333,16'd3002,16'd4252,-16'd449,16'd10123,16'd3066,16'd7117,-16'd1724,16'd617,-16'd5404,-16'd3563,16'd1940,-16'd441,16'd4654,16'd216,-16'd6150,-16'd5061,16'd1876,-16'd3736,-16'd756,-16'd5947,-16'd5542,-16'd952,-16'd5529,16'd1786};
dout[1023]={ 16'd1040,-16'd1981,-16'd1892,-16'd2086,16'd4023,-16'd6517,-16'd3556,-16'd2742,-16'd15615,16'd3504,16'd3753,16'd3353,-16'd3439,-16'd4894,16'd2523,-16'd4563,-16'd1186,16'd4925,16'd2745,-16'd10477,-16'd1298,16'd3863,16'd1318,-16'd2406,-16'd1750,-16'd696,-16'd8936,16'd8127,-16'd3892,-16'd4918,-16'd1532,-16'd5387,16'd207,16'd3852,-16'd776,16'd678};
dout[1024]={ 16'd6295,16'd1637,-16'd8718,-16'd6051,16'd666,-16'd4304,-16'd2700,16'd35,16'd267,16'd2376,16'd1112,-16'd2137,-16'd3083,16'd2354,-16'd2800,16'd4854,-16'd2130,-16'd7201,16'd1327,16'd408,-16'd1552,-16'd5995,-16'd7328,16'd11558,16'd4135,-16'd2908,-16'd8392,16'd6905,-16'd4756,-16'd358,16'd89,16'd3800,16'd2894,-16'd2604,-16'd5828,-16'd122};
dout[1025]={ 16'd1022,-16'd1229,-16'd5466,-16'd2583,16'd4477,-16'd4952,16'd2177,-16'd8239,-16'd2646,16'd2444,16'd3402,16'd7072,16'd1083,16'd4736,16'd3289,16'd2259,16'd569,-16'd3840,-16'd3428,-16'd1334,16'd3639,16'd4127,-16'd6556,-16'd2254,-16'd5722,-16'd3809,-16'd1880,16'd7235,16'd7627,-16'd8339,-16'd863,16'd5205,16'd6072,-16'd3513,-16'd876,16'd1610};
dout[1026]={ -16'd1115,-16'd2274,-16'd149,-16'd7494,-16'd2587,-16'd8764,-16'd324,-16'd6963,16'd4149,16'd641,16'd1771,-16'd4990,16'd505,-16'd4153,-16'd4102,16'd3989,-16'd8928,16'd5148,16'd5514,-16'd6941,-16'd8409,-16'd4555,16'd801,-16'd4644,-16'd5953,-16'd2471,-16'd4635,16'd1272,-16'd4388,-16'd6682,-16'd6136,-16'd6178,-16'd1158,16'd6581,-16'd1782,-16'd5267};
dout[1027]={ -16'd3136,16'd6162,16'd3707,-16'd7083,-16'd5846,16'd396,16'd1704,-16'd5773,16'd6676,-16'd5705,16'd3304,-16'd1376,16'd3187,16'd4738,-16'd391,16'd814,16'd1276,-16'd2170,16'd5903,16'd275,16'd293,-16'd7384,-16'd3410,16'd2080,16'd530,16'd1687,-16'd4650,-16'd1236,16'd4885,-16'd2406,-16'd760,16'd3181,-16'd4157,-16'd1497,16'd975,-16'd3596};
dout[1028]={ -16'd3081,16'd515,-16'd1232,-16'd10884,-16'd3220,-16'd540,-16'd5853,-16'd8606,16'd4446,16'd892,-16'd6698,16'd7137,-16'd3060,16'd1603,16'd4287,16'd6050,-16'd4867,16'd5069,-16'd2612,16'd7843,16'd3717,-16'd2152,-16'd287,-16'd6733,16'd7174,-16'd2042,16'd5639,16'd1795,16'd3199,16'd1282,16'd566,-16'd4628,16'd1881,16'd3152,16'd312,-16'd2098};
dout[1029]={ -16'd2631,16'd1544,16'd759,16'd2974,16'd2947,-16'd415,16'd2540,16'd1719,-16'd4366,-16'd2556,16'd3179,16'd5812,16'd181,16'd5319,-16'd2190,-16'd3301,-16'd6480,16'd6962,16'd2344,16'd6049,-16'd3269,16'd3720,16'd3849,-16'd2474,16'd1961,16'd2315,-16'd3805,-16'd7272,16'd6943,-16'd5886,-16'd4849,-16'd1484,16'd5338,-16'd993,-16'd1332,16'd88};
dout[1030]={ -16'd3780,-16'd9350,16'd1804,16'd7102,-16'd8113,-16'd5133,-16'd2451,16'd7990,16'd7178,-16'd2576,-16'd8193,16'd9479,16'd467,16'd6315,-16'd6447,16'd1375,-16'd2812,-16'd8526,16'd9212,16'd1034,16'd4119,-16'd2822,-16'd1220,16'd5506,16'd942,16'd3814,16'd4620,16'd910,-16'd3602,16'd2289,-16'd4958,-16'd2454,-16'd7173,-16'd2220,-16'd8700,-16'd7222};
dout[1031]={ -16'd5954,-16'd4326,-16'd2691,-16'd5056,-16'd6193,16'd6248,16'd3372,-16'd3591,16'd10343,-16'd11148,16'd2099,16'd6708,16'd6732,16'd5387,16'd4799,16'd7080,16'd3956,16'd1024,-16'd2587,-16'd28,16'd3394,-16'd594,16'd1246,-16'd2334,-16'd4286,16'd9495,16'd4023,-16'd1733,16'd4660,16'd5523,16'd2953,16'd2997,16'd2489,16'd4641,16'd1739,16'd6719};
dout[1032]={ -16'd7358,-16'd3106,16'd5481,16'd4915,-16'd9199,-16'd2701,16'd752,16'd529,-16'd6350,-16'd875,-16'd7607,16'd6126,-16'd5448,16'd6249,16'd3543,-16'd5328,-16'd7193,16'd3593,16'd1348,16'd2461,-16'd8221,-16'd1368,-16'd7129,-16'd3032,-16'd240,16'd784,-16'd1084,16'd3685,16'd2072,-16'd5647,-16'd2152,-16'd4684,-16'd9029,16'd7188,-16'd5458,-16'd3034};
dout[1033]={ -16'd7641,16'd7456,16'd1896,16'd108,-16'd4870,16'd6962,-16'd659,16'd2822,-16'd13042,-16'd6572,16'd514,16'd264,16'd4759,16'd2928,16'd6336,16'd2973,-16'd5290,16'd296,-16'd1962,-16'd9291,16'd4058,16'd3678,-16'd1303,-16'd771,-16'd4724,-16'd1869,-16'd3094,16'd4414,16'd4202,-16'd1282,-16'd384,-16'd6296,-16'd5047,16'd5182,-16'd5897,-16'd3766};
dout[1034]={ -16'd7516,16'd3916,-16'd4254,-16'd4574,16'd2025,16'd4797,-16'd3154,16'd6744,-16'd11546,-16'd2924,-16'd3792,16'd3177,16'd7048,16'd4037,16'd4126,16'd1678,16'd4548,-16'd11111,16'd1512,-16'd298,16'd3544,16'd275,-16'd3549,16'd2710,-16'd5570,-16'd3532,-16'd5659,16'd1537,-16'd5990,-16'd2153,16'd2000,16'd3614,-16'd8012,-16'd9618,-16'd582,-16'd5384};
dout[1035]={ -16'd8674,-16'd792,-16'd4,-16'd3585,16'd979,-16'd7673,-16'd5553,-16'd4612,-16'd1724,-16'd3872,16'd435,16'd4699,-16'd4328,-16'd3302,-16'd1987,16'd9268,-16'd7976,-16'd4557,-16'd4465,-16'd3803,16'd2365,16'd3563,16'd5265,16'd6648,16'd6215,16'd221,-16'd3353,16'd8021,-16'd1228,16'd2344,16'd1761,16'd1930,-16'd2772,-16'd3967,-16'd2126,16'd2902};
dout[1036]={ -16'd251,16'd1592,-16'd5321,-16'd997,16'd3162,-16'd1347,-16'd6071,16'd6413,16'd599,-16'd8644,16'd5505,16'd2979,16'd7028,16'd2470,-16'd2390,-16'd1717,16'd1770,-16'd8706,-16'd5459,16'd625,-16'd8474,16'd4884,-16'd7432,-16'd113,16'd6388,16'd1333,16'd2858,16'd6254,16'd1618,-16'd1105,-16'd3395,16'd5360,16'd5245,-16'd5870,-16'd4498,-16'd6461};
dout[1037]={ 16'd3588,16'd3723,-16'd6538,-16'd6557,16'd2725,-16'd2312,16'd2783,-16'd5058,-16'd2987,16'd3210,16'd4538,16'd2294,16'd2878,-16'd2721,-16'd4347,-16'd1174,16'd3715,16'd3859,16'd3923,16'd255,16'd600,-16'd2552,-16'd1804,16'd7189,16'd3788,16'd3915,16'd1169,16'd5435,16'd4420,-16'd4033,16'd4767,16'd8442,-16'd3561,16'd777,-16'd4665,16'd4213};
dout[1038]={ 16'd325,16'd1151,16'd1680,-16'd5790,16'd3051,-16'd8769,16'd7681,-16'd3833,-16'd4457,-16'd8810,-16'd6288,-16'd5704,-16'd232,16'd679,16'd3333,16'd1055,-16'd3493,16'd2711,-16'd5074,16'd2283,16'd4754,16'd1394,16'd5672,-16'd2069,16'd8376,16'd2256,16'd256,16'd1726,-16'd1458,16'd2015,-16'd3629,-16'd6946,16'd611,-16'd6435,-16'd2495,16'd5634};
dout[1039]={ 16'd5033,16'd2165,-16'd5630,-16'd3461,-16'd7838,-16'd11037,16'd5265,16'd2473,-16'd140,-16'd6040,16'd6992,-16'd2823,16'd6332,16'd4694,-16'd5049,16'd945,16'd2520,16'd6648,-16'd3731,16'd4187,16'd46,16'd3813,16'd6049,-16'd4731,-16'd2036,-16'd4216,-16'd4421,16'd3549,-16'd4357,-16'd3422,-16'd5880,-16'd1616,16'd5301,-16'd4249,16'd1496,-16'd3061};
dout[1040]={ 16'd4319,-16'd7055,-16'd9964,-16'd4857,-16'd4086,16'd7397,-16'd6170,16'd6400,16'd7034,-16'd95,-16'd4421,16'd10676,16'd4218,16'd428,-16'd5317,16'd10474,-16'd2565,16'd128,16'd2020,-16'd14654,-16'd5499,-16'd8293,-16'd3717,16'd3480,-16'd2471,16'd8568,-16'd3555,16'd8984,-16'd8795,16'd1236,16'd4411,16'd5076,16'd4795,-16'd11475,16'd3943,-16'd2101};
dout[1041]={ -16'd2843,-16'd1650,16'd7975,16'd8549,16'd5461,16'd1124,-16'd340,16'd2087,16'd5357,-16'd8575,16'd4708,-16'd3155,16'd4238,-16'd8543,16'd3962,16'd5806,16'd3271,16'd2519,-16'd2015,-16'd4343,-16'd2860,-16'd4125,-16'd4367,-16'd5465,16'd6293,-16'd1406,-16'd5913,-16'd2667,16'd6257,16'd885,16'd1459,16'd2541,-16'd6697,16'd2052,16'd1915,16'd3057};
dout[1042]={ 16'd3773,16'd6366,16'd7721,-16'd1497,-16'd6670,16'd3645,16'd6721,16'd3359,16'd2687,16'd1860,16'd369,-16'd5654,16'd6448,16'd5907,-16'd6549,-16'd4386,16'd2215,16'd5831,-16'd149,-16'd7276,16'd5657,-16'd5463,-16'd4029,-16'd7425,16'd1139,-16'd2488,-16'd7634,16'd4144,16'd4500,16'd6272,-16'd2289,16'd2781,16'd1388,-16'd4857,16'd7771,16'd6537};
dout[1043]={ -16'd656,16'd136,16'd4031,16'd9172,16'd259,-16'd31,-16'd2646,16'd371,-16'd15092,-16'd8553,-16'd4109,-16'd1660,16'd6016,16'd1778,-16'd2055,-16'd4122,16'd3839,16'd3934,-16'd7130,-16'd9948,-16'd2277,-16'd7604,-16'd3733,16'd1066,-16'd3379,-16'd3483,-16'd3694,16'd2756,-16'd1701,16'd6927,16'd3677,-16'd887,16'd4006,-16'd5696,16'd5159,16'd2992};
dout[1044]={ -16'd3244,-16'd4950,16'd2127,-16'd3637,-16'd1150,16'd6217,-16'd218,16'd4501,-16'd2974,-16'd1532,-16'd6897,16'd8373,-16'd4147,-16'd675,-16'd6825,16'd6912,-16'd5439,-16'd4560,-16'd6086,-16'd6400,-16'd7755,16'd2287,-16'd3286,16'd7787,16'd3462,16'd1501,-16'd123,16'd4021,16'd7040,16'd1353,16'd3668,16'd7666,-16'd3970,-16'd5254,-16'd2507,-16'd7752};
dout[1045]={ -16'd426,16'd4565,-16'd7634,16'd608,16'd5142,16'd586,-16'd7655,16'd2827,-16'd4142,-16'd4278,-16'd8447,-16'd1294,16'd5551,16'd2139,16'd4741,16'd7707,16'd6741,-16'd1864,16'd8409,-16'd2698,16'd2910,16'd4275,16'd4515,-16'd2887,-16'd2315,-16'd155,-16'd4412,-16'd1901,-16'd3148,16'd3015,16'd111,-16'd4514,-16'd8254,16'd2832,16'd4719,16'd5924};
dout[1046]={ -16'd2343,16'd6396,-16'd1291,-16'd8230,-16'd6124,16'd1598,16'd1621,16'd2604,-16'd6157,-16'd2696,-16'd6400,16'd6026,-16'd1000,16'd4877,-16'd838,16'd2205,-16'd75,-16'd6656,-16'd6500,-16'd235,-16'd1875,-16'd344,16'd5399,16'd958,16'd7245,-16'd2613,16'd353,-16'd1863,16'd6276,-16'd8150,16'd4762,16'd1239,16'd1501,-16'd7223,16'd3247,16'd2056};
dout[1047]={ 16'd2497,-16'd6264,16'd357,-16'd6583,-16'd8106,16'd1224,16'd1453,16'd1697,-16'd3777,16'd7558,-16'd2094,-16'd1912,16'd7455,-16'd7392,16'd1077,16'd946,16'd5434,-16'd3424,16'd4048,16'd730,16'd2211,16'd2290,-16'd3861,-16'd5871,-16'd1775,16'd5461,-16'd5604,-16'd3655,16'd5931,-16'd7244,16'd4064,-16'd4423,16'd976,16'd831,-16'd1811,16'd2838};
dout[1048]={ -16'd3773,-16'd4831,-16'd8625,-16'd4104,-16'd9336,-16'd1159,16'd2887,-16'd482,16'd6,-16'd4879,-16'd4007,16'd6933,-16'd6355,16'd5636,16'd263,16'd1277,16'd3023,-16'd4055,-16'd1425,-16'd5406,16'd5591,16'd5126,16'd3805,16'd5888,-16'd940,16'd4677,-16'd2569,16'd749,16'd4848,-16'd154,16'd176,16'd6651,-16'd6278,16'd343,-16'd8157,-16'd5496};
dout[1049]={ -16'd5828,16'd492,-16'd1867,16'd4413,16'd2740,16'd1175,16'd5111,-16'd6402,-16'd141,-16'd1236,-16'd5644,16'd2148,16'd6164,-16'd4415,-16'd2900,-16'd598,-16'd5702,-16'd4325,16'd1697,-16'd2557,-16'd3059,-16'd4315,-16'd5809,16'd5979,-16'd4701,16'd4957,16'd4361,-16'd1366,-16'd1556,-16'd3824,16'd6432,16'd4970,-16'd7373,16'd1252,16'd1828,16'd2124};
dout[1050]={ -16'd2885,16'd1453,-16'd8030,16'd1363,-16'd960,-16'd5232,-16'd1473,16'd6884,16'd6969,-16'd4052,-16'd9562,16'd1864,16'd12036,16'd2913,-16'd4557,16'd10585,-16'd1031,-16'd8368,-16'd557,-16'd16489,-16'd5978,16'd3989,-16'd9594,16'd11030,16'd2926,16'd3894,-16'd6969,16'd7678,-16'd10424,16'd43,16'd6284,16'd6380,16'd2222,-16'd6053,16'd6223,-16'd2673};
dout[1051]={ -16'd3146,-16'd8552,16'd1270,16'd4647,-16'd1184,-16'd7487,-16'd3058,16'd1190,16'd9940,-16'd8113,-16'd470,-16'd74,-16'd408,-16'd4828,-16'd5199,16'd1681,16'd5870,16'd3361,16'd4642,-16'd3136,-16'd7657,16'd4529,-16'd3222,-16'd2422,16'd3042,16'd3322,-16'd3980,-16'd3781,-16'd1488,16'd2383,16'd6890,16'd1619,-16'd8060,-16'd2813,-16'd314,-16'd2516};
dout[1052]={ -16'd1319,-16'd5093,16'd3788,16'd2525,-16'd5320,-16'd8372,-16'd2335,16'd2275,16'd7449,16'd1599,-16'd4374,16'd1007,16'd325,-16'd3220,-16'd3664,-16'd3933,16'd7098,-16'd3686,16'd5718,-16'd8185,16'd5,-16'd7226,16'd1463,-16'd4121,16'd4953,-16'd7062,-16'd7179,16'd8058,16'd2345,-16'd2562,16'd2675,16'd499,-16'd7399,-16'd742,-16'd344,16'd2815};
dout[1053]={ -16'd495,16'd3412,-16'd1714,-16'd2474,-16'd4430,-16'd8646,-16'd657,16'd7767,-16'd3018,16'd1321,-16'd7455,-16'd6131,-16'd4583,-16'd5986,-16'd25,16'd8534,-16'd184,-16'd6139,16'd2475,16'd3055,16'd3984,-16'd3936,16'd1742,16'd5160,16'd4732,16'd812,-16'd6260,-16'd383,-16'd735,-16'd5023,16'd6838,16'd5633,16'd4394,16'd3723,16'd4564,16'd4131};
dout[1054]={ -16'd5971,-16'd2413,-16'd2178,16'd6945,16'd2610,-16'd8498,16'd3909,16'd1915,-16'd643,16'd1735,-16'd9074,-16'd3912,16'd2345,16'd8659,-16'd857,16'd2407,16'd5332,-16'd6215,-16'd3071,16'd3070,16'd3748,-16'd6106,-16'd6848,-16'd4674,-16'd4848,16'd6863,16'd3882,16'd4099,-16'd6501,16'd3952,16'd6005,16'd5239,-16'd8339,-16'd2055,16'd1603,16'd4524};
dout[1055]={ -16'd7917,16'd1302,-16'd7043,-16'd1828,16'd829,-16'd2278,16'd3051,-16'd1479,16'd6316,16'd814,-16'd9379,16'd5294,16'd5513,16'd2408,16'd4420,-16'd205,-16'd1402,-16'd189,-16'd5709,16'd216,-16'd4433,16'd3606,-16'd4010,16'd5479,16'd7435,-16'd855,-16'd2494,16'd4465,-16'd2597,16'd2206,16'd1601,16'd4823,-16'd7889,16'd4822,16'd985,-16'd6393};
dout[1056]={ -16'd4210,-16'd3523,16'd4986,-16'd1232,16'd1395,-16'd8562,-16'd6867,16'd3514,16'd5362,-16'd1187,-16'd5178,-16'd1559,-16'd654,16'd4099,-16'd1018,16'd5293,-16'd1803,-16'd5755,16'd2881,16'd2405,-16'd8095,-16'd810,-16'd1899,-16'd17,16'd498,16'd1919,16'd3302,16'd727,16'd4361,16'd4801,-16'd6652,16'd901,16'd1227,-16'd6388,-16'd1904,16'd5860};
dout[1057]={ 16'd1845,-16'd1000,-16'd1529,-16'd2315,16'd2465,-16'd2374,-16'd48,16'd158,-16'd7658,16'd8730,16'd2602,-16'd65,-16'd1433,16'd6961,-16'd6251,16'd4183,-16'd1476,-16'd7048,-16'd2345,-16'd4862,-16'd3038,16'd2791,16'd797,16'd2744,-16'd5944,-16'd4115,16'd1469,16'd2646,-16'd5010,-16'd981,16'd19,-16'd4480,-16'd8817,-16'd6735,16'd3238,16'd3627};
dout[1058]={ -16'd5231,16'd4763,-16'd1855,16'd354,16'd4992,-16'd4302,-16'd602,16'd3522,-16'd6485,16'd7303,-16'd327,-16'd5941,16'd4959,-16'd705,-16'd9872,-16'd325,16'd540,16'd3199,16'd3102,-16'd1522,-16'd3643,16'd3719,16'd3472,-16'd5159,-16'd5073,-16'd2449,-16'd2853,-16'd4853,16'd537,16'd4061,16'd2963,-16'd4471,-16'd7591,16'd1288,-16'd539,-16'd2719};
dout[1059]={ 16'd1192,-16'd6205,-16'd3208,-16'd5474,-16'd2382,-16'd11461,16'd7593,-16'd2074,-16'd2413,16'd6333,16'd3717,16'd1604,-16'd5029,16'd1081,-16'd7094,-16'd6999,16'd2225,16'd6582,16'd2054,16'd6271,-16'd1574,-16'd7212,16'd1860,16'd6921,16'd8227,16'd1894,16'd5129,-16'd1125,-16'd4598,-16'd7603,16'd2647,-16'd2312,-16'd4224,-16'd8566,16'd3316,-16'd278};
dout[1060]={ 16'd5826,-16'd1509,16'd3153,16'd314,-16'd1165,-16'd1934,-16'd8956,16'd1481,16'd711,16'd1309,-16'd8281,-16'd3165,16'd13869,-16'd598,16'd520,16'd1124,16'd4129,-16'd2751,16'd8332,-16'd5798,16'd27,-16'd562,-16'd8502,16'd12514,16'd1956,-16'd4170,16'd797,16'd8920,16'd3343,16'd247,-16'd4474,16'd5946,-16'd1731,-16'd476,16'd590,-16'd4991};
dout[1061]={ 16'd6205,-16'd4259,16'd5619,16'd3452,-16'd1832,-16'd7333,-16'd1568,16'd2759,16'd6912,16'd3181,16'd3894,-16'd982,16'd5316,-16'd10708,16'd3340,16'd3236,16'd7111,-16'd8344,16'd3489,-16'd6201,-16'd9352,-16'd8346,16'd3110,-16'd791,16'd3545,16'd6801,-16'd4013,-16'd4656,-16'd5038,-16'd7253,16'd621,16'd1862,-16'd3041,-16'd8471,-16'd760,16'd3099};
dout[1062]={ 16'd5302,16'd6432,16'd10184,16'd2026,16'd2811,16'd600,16'd197,-16'd2365,-16'd1194,-16'd5866,16'd945,-16'd5020,-16'd5424,-16'd4878,-16'd8834,-16'd100,-16'd4403,-16'd3182,-16'd8703,16'd3690,16'd3787,16'd3030,16'd6405,-16'd2910,16'd2546,-16'd2305,16'd1927,16'd3534,-16'd8285,-16'd7048,-16'd6118,-16'd7302,-16'd8256,-16'd732,-16'd6178,-16'd4116};
dout[1063]={ 16'd5865,-16'd38,16'd1546,16'd4143,-16'd4716,16'd1074,-16'd5339,16'd4029,-16'd9855,16'd4957,-16'd5664,-16'd7507,-16'd3726,16'd6449,-16'd4943,16'd1899,16'd180,-16'd8378,-16'd5853,16'd1410,-16'd3879,16'd2713,16'd1181,-16'd7281,16'd5893,-16'd3449,-16'd6041,16'd5016,16'd2982,-16'd1380,16'd5076,16'd3110,-16'd2959,-16'd495,-16'd2099,-16'd9362};
dout[1064]={ -16'd4693,-16'd5485,-16'd3401,16'd4205,16'd1753,16'd342,-16'd2560,-16'd2889,-16'd8329,-16'd6757,16'd3088,-16'd624,-16'd1864,-16'd514,-16'd3346,-16'd1121,16'd3596,-16'd9788,-16'd2535,-16'd933,-16'd5070,16'd4405,-16'd2797,16'd4836,-16'd2088,16'd2169,16'd5735,-16'd1989,-16'd5662,16'd2249,16'd535,16'd4749,-16'd4295,-16'd2343,-16'd3826,-16'd1433};
dout[1065]={ 16'd5484,16'd1081,16'd1008,16'd2928,-16'd6346,-16'd5539,16'd2455,16'd665,-16'd3031,-16'd5152,-16'd4606,16'd4282,16'd1872,-16'd1424,-16'd1719,16'd1424,16'd726,-16'd3692,16'd2853,-16'd5766,16'd5028,16'd407,-16'd5487,-16'd192,-16'd3768,16'd5894,16'd6893,16'd6216,16'd4525,-16'd6905,16'd5307,-16'd4106,-16'd3564,-16'd4970,-16'd8381,-16'd4732};
dout[1066]={ -16'd6048,-16'd5951,16'd98,16'd2694,16'd2856,-16'd5375,-16'd6933,16'd4745,16'd3003,16'd7406,-16'd387,16'd2267,-16'd2865,16'd3106,16'd3625,16'd2134,-16'd2963,-16'd9053,16'd5700,16'd2022,-16'd4418,16'd1076,-16'd5210,16'd2416,16'd908,-16'd3560,-16'd714,-16'd2640,-16'd5155,-16'd5854,-16'd5185,-16'd5188,-16'd3946,16'd4638,-16'd7182,-16'd5670};
dout[1067]={ 16'd1124,-16'd4492,16'd1696,-16'd648,-16'd6731,16'd2764,-16'd1694,16'd4184,-16'd2545,-16'd596,16'd3471,16'd38,16'd6786,-16'd2279,-16'd9003,16'd528,16'd2230,-16'd5621,16'd4115,16'd1452,16'd1894,16'd2657,16'd5625,16'd5851,16'd164,16'd566,-16'd5544,-16'd605,16'd3276,16'd5023,16'd2807,-16'd1018,16'd1985,-16'd9128,16'd1892,-16'd3946};
dout[1068]={ -16'd876,-16'd1490,16'd486,-16'd1751,-16'd4798,-16'd3644,-16'd2096,16'd2551,16'd8338,-16'd2217,-16'd3539,16'd1907,16'd4666,-16'd7110,16'd1744,-16'd50,-16'd6179,-16'd4680,16'd4170,16'd2993,16'd495,16'd5862,16'd4452,16'd1078,-16'd2203,-16'd5463,-16'd674,-16'd3233,16'd1774,-16'd3752,16'd1791,16'd2944,-16'd8242,-16'd2208,16'd6913,-16'd4122};
dout[1069]={ -16'd6573,16'd178,-16'd399,-16'd3559,-16'd2057,16'd2272,16'd4687,16'd1340,16'd4438,16'd5354,16'd460,16'd2046,-16'd5580,16'd4327,-16'd8290,16'd6490,16'd2874,16'd2624,-16'd5144,-16'd313,16'd1206,16'd4271,-16'd4177,16'd7141,16'd221,16'd8489,16'd824,16'd562,16'd7693,16'd369,16'd1535,-16'd2012,-16'd255,-16'd3587,-16'd2524,-16'd5011};
dout[1070]={ -16'd888,-16'd3640,-16'd6362,16'd455,16'd1384,16'd5761,-16'd5140,16'd9616,16'd9123,16'd4085,-16'd7034,-16'd5020,16'd474,-16'd3362,16'd6395,-16'd1669,-16'd3716,-16'd9822,16'd1994,16'd1825,16'd6770,16'd3325,-16'd10523,16'd9911,16'd1235,-16'd8477,16'd5438,16'd3714,-16'd703,16'd5600,16'd6696,16'd1802,-16'd2567,16'd4121,-16'd5918,16'd5504};
dout[1071]={ -16'd5163,16'd1597,16'd804,16'd745,16'd2131,16'd1604,16'd6173,16'd6439,16'd8746,-16'd1477,-16'd8568,16'd2514,-16'd8046,-16'd947,-16'd5179,16'd8243,16'd1764,16'd3195,-16'd2336,16'd5328,16'd331,-16'd1953,-16'd4250,-16'd4056,-16'd1033,-16'd5448,-16'd1221,16'd6360,16'd1322,-16'd854,-16'd6200,16'd2775,16'd3349,-16'd4031,-16'd7894,-16'd1912};
dout[1072]={ 16'd5428,16'd4564,16'd3035,16'd1053,-16'd6961,-16'd170,16'd3486,-16'd2114,16'd4321,16'd4184,16'd861,16'd4051,-16'd8607,16'd836,16'd2609,16'd1700,-16'd6282,-16'd6128,-16'd7863,16'd3785,-16'd5045,16'd4184,-16'd3832,-16'd6391,16'd5996,16'd2916,-16'd6954,-16'd404,-16'd7430,-16'd800,16'd1490,-16'd8014,-16'd3393,16'd2235,-16'd751,16'd2663};
dout[1073]={ 16'd4624,16'd1007,16'd9439,16'd5010,-16'd4489,16'd508,-16'd3010,16'd2128,-16'd2836,-16'd3578,-16'd5284,16'd2043,16'd1624,-16'd1579,16'd1051,16'd376,-16'd5207,-16'd6814,-16'd9206,-16'd1899,-16'd4147,-16'd2523,16'd5140,16'd1037,-16'd2774,-16'd140,-16'd6561,-16'd4154,-16'd7080,16'd646,16'd6902,16'd7624,16'd2614,-16'd3033,-16'd5187,16'd3321};
dout[1074]={ -16'd1815,-16'd8025,16'd8262,-16'd5575,-16'd2621,16'd4671,-16'd7510,16'd8501,-16'd2924,16'd6171,16'd4177,-16'd3661,16'd3067,16'd4179,16'd6053,16'd3341,16'd3673,-16'd3815,16'd2148,16'd1470,-16'd576,16'd1325,-16'd7303,16'd4811,16'd6989,-16'd3462,-16'd4107,-16'd7584,16'd2514,-16'd3379,16'd4951,16'd2061,16'd57,-16'd1824,16'd132,16'd3368};
dout[1075]={ 16'd2651,16'd1234,-16'd2814,-16'd2419,-16'd2342,16'd2741,16'd3423,16'd6590,-16'd138,-16'd1878,-16'd2779,-16'd2631,-16'd2575,-16'd794,-16'd8430,-16'd6764,16'd4733,16'd2340,-16'd495,16'd7353,-16'd2913,-16'd4189,-16'd6870,16'd1525,-16'd4810,-16'd2196,-16'd3475,-16'd4309,-16'd3732,16'd7576,16'd4569,-16'd8095,-16'd3350,-16'd5699,-16'd1670,16'd3562};
dout[1076]={ 16'd650,-16'd1472,-16'd4974,16'd4685,-16'd892,16'd1616,-16'd1151,16'd2688,16'd6359,-16'd546,16'd4638,16'd2126,16'd2541,-16'd1282,-16'd7892,-16'd3483,16'd4416,-16'd1104,16'd2992,16'd4191,16'd7976,16'd6145,-16'd2348,-16'd3737,16'd6202,16'd6008,16'd6847,-16'd3101,16'd4401,-16'd3450,-16'd3663,16'd3234,-16'd6764,-16'd3922,-16'd2967,-16'd7178};
dout[1077]={ -16'd3955,16'd3479,-16'd546,16'd2842,16'd125,16'd2224,-16'd2925,16'd2799,-16'd4824,16'd4932,16'd68,-16'd5915,-16'd1506,16'd4998,16'd198,16'd537,16'd1589,-16'd9864,16'd311,-16'd5249,16'd633,-16'd3729,-16'd7353,-16'd1753,-16'd751,-16'd4084,16'd6999,16'd2598,-16'd4537,16'd2922,-16'd5207,-16'd552,-16'd2983,16'd3809,-16'd5986,16'd3597};
dout[1078]={ -16'd4994,-16'd4014,16'd1883,-16'd2165,16'd2228,-16'd8091,16'd1564,-16'd3613,16'd7534,16'd3785,16'd1949,-16'd361,-16'd8343,-16'd8054,16'd4144,-16'd2328,-16'd6808,16'd3260,16'd3874,-16'd4771,16'd3160,16'd8657,16'd946,16'd4918,-16'd6454,16'd2458,-16'd1511,-16'd2569,16'd6519,16'd3685,16'd6165,16'd131,-16'd4230,16'd2734,16'd5464,16'd792};
dout[1079]={ 16'd2488,-16'd4344,-16'd1524,16'd1170,16'd4099,-16'd5143,-16'd5752,16'd4766,16'd3418,16'd425,-16'd2290,-16'd8422,16'd1306,-16'd4733,-16'd112,-16'd5357,-16'd1511,-16'd5416,16'd1393,16'd4569,16'd1437,-16'd4256,-16'd6364,16'd4644,-16'd6707,-16'd796,16'd8682,-16'd332,-16'd2400,-16'd3083,16'd4816,16'd3212,16'd4424,-16'd3413,-16'd6377,16'd1021};
dout[1080]={ 16'd400,-16'd10847,-16'd5583,16'd1289,-16'd1585,16'd5318,16'd5958,16'd3194,16'd5615,-16'd2601,16'd415,-16'd1268,16'd4464,-16'd4292,-16'd759,-16'd3646,16'd5997,16'd4488,-16'd679,-16'd866,16'd5183,16'd7005,-16'd4888,16'd12344,-16'd4970,16'd2965,16'd1105,-16'd701,16'd898,16'd347,-16'd1021,16'd2885,16'd2351,-16'd2082,16'd4352,16'd787};
dout[1081]={ 16'd4912,-16'd4528,-16'd8117,-16'd1244,-16'd2690,16'd1798,16'd4261,16'd5266,-16'd382,-16'd1103,-16'd3778,16'd969,-16'd6971,16'd4283,16'd4687,-16'd2479,16'd5508,-16'd482,-16'd4564,-16'd4352,16'd6611,16'd6007,-16'd9135,16'd3926,16'd8022,-16'd1290,-16'd5427,16'd1863,-16'd8551,-16'd4403,-16'd4717,16'd6527,-16'd8871,16'd675,-16'd701,-16'd6173};
dout[1082]={ -16'd4079,-16'd2360,-16'd3661,-16'd5148,16'd6461,-16'd2409,16'd4364,-16'd7212,-16'd2828,-16'd372,-16'd1910,16'd269,-16'd11427,16'd1202,-16'd4762,16'd4313,-16'd1595,16'd6019,16'd5745,16'd3889,16'd495,16'd1069,16'd5059,16'd4011,16'd8965,16'd3502,16'd3495,-16'd3677,-16'd9808,16'd2191,16'd3776,-16'd5952,-16'd5084,16'd4648,-16'd9154,16'd1184};
dout[1083]={ 16'd7029,-16'd3149,16'd7427,-16'd4746,-16'd5272,16'd4043,16'd632,-16'd5248,16'd4566,16'd1678,-16'd1510,-16'd8651,-16'd2522,16'd481,16'd2863,16'd6429,16'd4573,16'd1592,-16'd5375,-16'd1866,-16'd5663,16'd3767,16'd6814,16'd1241,16'd317,-16'd1536,-16'd3508,16'd1794,-16'd3662,-16'd3787,-16'd2261,-16'd3542,16'd991,-16'd939,16'd4203,-16'd337};
dout[1084]={ 16'd5970,-16'd3201,16'd2358,-16'd4517,16'd5537,-16'd1519,16'd3995,-16'd617,-16'd8328,-16'd3723,-16'd4808,16'd1090,-16'd1503,16'd346,-16'd7183,-16'd6594,-16'd6726,16'd3903,-16'd412,16'd563,16'd287,16'd8210,-16'd3167,16'd1322,16'd3073,16'd5661,16'd6015,-16'd9123,-16'd3481,-16'd273,16'd3423,16'd3372,-16'd2288,-16'd2733,-16'd5697,-16'd6749};
dout[1085]={ 16'd2362,16'd4306,-16'd197,16'd8202,16'd1279,16'd5955,-16'd4836,16'd1012,16'd7247,16'd1472,-16'd4809,-16'd1290,-16'd5303,-16'd1722,-16'd6675,-16'd7975,-16'd3011,-16'd3397,-16'd1188,-16'd3684,16'd5530,-16'd4520,16'd4071,-16'd3759,16'd2038,16'd2025,-16'd6114,16'd4545,-16'd6526,16'd8222,-16'd847,-16'd9004,16'd3428,16'd3172,16'd3527,-16'd4814};
dout[1086]={ 16'd3914,16'd491,16'd6187,16'd7724,-16'd6813,-16'd1495,16'd5542,-16'd5614,-16'd4603,16'd982,16'd1347,-16'd383,-16'd8474,-16'd7647,-16'd4412,-16'd269,16'd7052,-16'd3776,-16'd1702,16'd1747,-16'd4618,16'd2011,-16'd7125,-16'd3479,16'd1622,16'd2112,16'd5881,16'd2548,-16'd1712,16'd7221,16'd3931,-16'd9397,16'd365,16'd3400,16'd1828,16'd1440};
dout[1087]={ -16'd1487,16'd1503,-16'd6626,16'd4671,-16'd596,16'd3241,-16'd1225,-16'd666,-16'd2668,-16'd7270,16'd2765,16'd5351,-16'd9643,-16'd392,-16'd3464,16'd953,-16'd7272,-16'd1917,16'd450,-16'd2312,16'd4135,-16'd1464,-16'd6112,16'd2966,-16'd1232,16'd3775,-16'd2601,16'd5941,16'd597,-16'd2890,16'd3614,-16'd4207,16'd4963,-16'd9406,16'd3830,-16'd6185};
dout[1088]={ -16'd4639,-16'd6408,16'd6053,16'd4550,-16'd5660,16'd3559,16'd5491,-16'd1396,-16'd2459,-16'd564,-16'd5171,-16'd908,-16'd5661,-16'd7337,16'd989,-16'd2717,16'd1256,-16'd2783,-16'd3831,16'd4986,-16'd5866,16'd1061,16'd4428,-16'd393,16'd3110,-16'd1180,16'd3677,16'd2903,16'd3915,-16'd3207,16'd1654,16'd1874,-16'd6765,-16'd4323,-16'd9899,-16'd1066};
dout[1089]={ 16'd3658,16'd293,16'd7358,-16'd4399,-16'd7267,-16'd964,16'd6500,-16'd2288,-16'd3182,-16'd4415,-16'd3004,16'd2156,-16'd9023,-16'd3704,-16'd6480,16'd4296,16'd3174,-16'd1912,-16'd4958,16'd909,16'd7955,16'd2879,-16'd4356,-16'd5546,16'd534,16'd793,16'd7118,16'd3330,16'd5531,-16'd2857,-16'd6631,16'd5966,-16'd2019,-16'd4077,-16'd6080,-16'd1680};
dout[1090]={ -16'd3529,16'd436,-16'd7013,16'd1946,-16'd3214,16'd1618,16'd5216,16'd1782,16'd5145,16'd5129,-16'd1526,-16'd2168,16'd2661,-16'd4284,-16'd6135,-16'd15163,16'd887,-16'd3378,16'd963,-16'd9782,16'd5422,16'd3489,-16'd5645,16'd12625,-16'd6200,-16'd6338,16'd1149,16'd7245,-16'd5454,16'd3120,16'd3336,16'd611,-16'd8421,16'd7220,16'd2857,16'd6929};
dout[1091]={ -16'd7621,16'd5563,16'd0,-16'd3134,16'd156,-16'd7542,-16'd3195,16'd5670,-16'd5088,-16'd8635,-16'd7253,16'd6479,16'd2008,-16'd6969,16'd1045,16'd4776,-16'd5656,-16'd3784,16'd4126,16'd3562,-16'd1946,16'd4059,16'd2883,-16'd2277,16'd647,16'd1487,-16'd8225,-16'd5161,16'd1871,16'd1163,16'd7378,16'd2347,-16'd6138,16'd7789,-16'd8409,-16'd8090};
dout[1092]={ -16'd6106,-16'd4404,-16'd7486,-16'd2869,16'd7698,-16'd1983,-16'd810,-16'd10501,16'd1191,-16'd6242,-16'd3095,16'd1042,-16'd1853,16'd5753,-16'd4930,-16'd4255,-16'd4059,-16'd5593,-16'd2400,16'd4640,16'd6105,16'd2093,16'd1468,16'd1685,-16'd991,-16'd8450,-16'd3450,16'd2300,-16'd7331,16'd5677,16'd1888,-16'd3452,-16'd7791,16'd9358,-16'd9131,16'd369};
dout[1093]={ -16'd661,16'd6247,16'd9189,16'd5643,-16'd5346,16'd3605,-16'd1532,-16'd9081,-16'd7211,16'd5383,-16'd5414,-16'd8036,-16'd5861,-16'd581,-16'd5754,-16'd6228,16'd7284,16'd217,-16'd1780,16'd5029,-16'd3770,16'd4226,16'd6507,16'd2102,16'd6580,16'd5782,-16'd691,-16'd839,-16'd4756,-16'd10918,16'd4959,16'd2186,-16'd1758,16'd3953,-16'd8162,-16'd2314};
dout[1094]={ 16'd5160,-16'd9422,16'd1013,-16'd4900,16'd1873,-16'd58,16'd1774,-16'd4197,-16'd4696,16'd6191,-16'd5886,16'd6155,-16'd3989,-16'd5628,-16'd1734,-16'd7747,16'd683,-16'd5450,16'd5752,16'd6939,-16'd3378,16'd1478,-16'd7275,16'd3532,-16'd690,16'd9170,16'd4664,-16'd4129,16'd4672,-16'd10595,-16'd5330,16'd1361,16'd4047,16'd2611,16'd4418,16'd5091};
dout[1095]={ 16'd2389,16'd3130,-16'd842,-16'd3698,-16'd751,-16'd6517,-16'd1327,-16'd2290,16'd1385,16'd4298,16'd2689,16'd4448,-16'd8098,16'd2250,16'd4055,16'd2860,-16'd4222,-16'd4400,-16'd5004,16'd3546,16'd3123,-16'd6898,-16'd6370,16'd2161,16'd8575,16'd122,16'd5654,16'd2539,-16'd8430,16'd59,16'd1838,16'd3133,-16'd4411,-16'd786,16'd1453,-16'd192};
dout[1096]={ 16'd4890,-16'd539,16'd3651,-16'd5347,16'd972,-16'd1011,-16'd2803,-16'd556,-16'd3643,-16'd1321,16'd4816,-16'd611,-16'd8505,-16'd4632,-16'd3961,-16'd6083,-16'd664,-16'd2389,16'd951,-16'd5164,16'd1244,-16'd4278,-16'd4972,16'd1463,-16'd4636,-16'd409,16'd4203,16'd858,-16'd3840,-16'd3137,-16'd1439,-16'd6309,-16'd628,16'd2316,-16'd879,-16'd5141};
dout[1097]={ 16'd1140,16'd2616,-16'd1282,16'd5038,-16'd2600,-16'd8072,16'd2942,16'd4161,16'd405,-16'd3574,-16'd3295,-16'd5266,-16'd7032,16'd7642,-16'd81,-16'd5737,-16'd6454,-16'd805,16'd3414,16'd7118,-16'd4513,-16'd6874,-16'd3078,-16'd2743,-16'd667,16'd147,16'd2873,-16'd4222,16'd2119,-16'd1141,16'd5216,-16'd7044,-16'd6763,-16'd2505,16'd1529,16'd2543};
dout[1098]={ -16'd1555,16'd2613,16'd2458,16'd5571,-16'd3245,16'd2220,-16'd2395,16'd1700,16'd2999,-16'd2360,-16'd7721,-16'd6191,16'd2666,16'd6573,-16'd493,16'd1118,-16'd6923,-16'd2694,16'd5976,-16'd5735,-16'd7969,16'd1709,16'd5815,16'd7248,-16'd3237,16'd949,-16'd7017,16'd3004,16'd5048,-16'd3475,-16'd1497,16'd1677,-16'd553,-16'd2740,-16'd3957,16'd2614};
dout[1099]={ -16'd308,-16'd2062,-16'd765,-16'd3915,-16'd8621,-16'd3444,16'd5071,-16'd1332,-16'd4927,16'd883,-16'd3416,16'd2577,16'd2487,-16'd7579,-16'd4903,16'd5081,-16'd5326,-16'd6450,-16'd4775,-16'd1543,-16'd1006,16'd3884,-16'd7132,16'd5755,16'd6515,16'd2612,-16'd2414,16'd206,16'd3728,-16'd5568,16'd430,16'd6167,-16'd971,16'd2025,-16'd7758,-16'd4008};
dout[1100]={ 16'd836,16'd641,-16'd8691,16'd3494,-16'd1841,16'd347,-16'd361,16'd7,-16'd6325,-16'd4722,-16'd6768,16'd247,-16'd186,-16'd356,16'd4283,-16'd15853,-16'd2914,-16'd5645,16'd5330,16'd3509,-16'd6921,16'd3516,-16'd5187,16'd10394,-16'd10149,-16'd8766,16'd5426,16'd2021,16'd1142,-16'd2144,16'd6717,-16'd3730,-16'd4316,16'd3037,16'd3482,-16'd2734};
dout[1101]={ -16'd1622,16'd6979,-16'd4253,-16'd9684,-16'd1092,16'd4198,-16'd7062,-16'd6481,16'd1962,-16'd1749,-16'd1714,-16'd1290,-16'd3313,16'd3967,16'd927,-16'd3656,-16'd270,-16'd6709,16'd486,-16'd1256,16'd4651,16'd5230,-16'd4652,16'd510,-16'd8787,-16'd4628,16'd6356,-16'd2350,-16'd3505,16'd1181,-16'd1434,-16'd6628,-16'd8003,16'd9035,-16'd647,16'd321};
dout[1102]={ -16'd8663,16'd2644,-16'd2108,-16'd2390,16'd5793,-16'd2666,16'd3903,-16'd10989,16'd958,-16'd10175,16'd2400,16'd6976,16'd3548,-16'd437,16'd4837,-16'd1570,-16'd3272,16'd4941,-16'd6996,-16'd206,-16'd1624,-16'd7260,-16'd2037,-16'd3111,16'd6914,-16'd6544,16'd704,16'd2038,16'd1911,-16'd9127,16'd9900,-16'd8238,16'd2961,16'd6176,16'd2524,-16'd1278};
dout[1103]={ -16'd8099,-16'd6053,-16'd5729,-16'd8074,16'd5617,16'd3978,-16'd940,-16'd9678,16'd2279,-16'd8667,-16'd8458,16'd3349,16'd3302,-16'd7295,16'd4192,16'd421,-16'd6331,16'd990,-16'd7945,16'd1915,-16'd1076,-16'd4040,-16'd2898,-16'd1062,16'd6181,-16'd3995,16'd81,16'd3719,16'd3500,-16'd7369,16'd6703,-16'd4802,-16'd3327,-16'd6602,16'd711,16'd5392};
dout[1104]={ -16'd5069,-16'd10089,16'd4683,16'd2778,-16'd4023,16'd3251,-16'd156,16'd3757,16'd2530,16'd4179,16'd5698,16'd249,-16'd1720,-16'd5429,-16'd8624,-16'd2404,16'd666,-16'd3507,-16'd2634,-16'd5439,-16'd5584,16'd2148,16'd294,-16'd4042,16'd2746,16'd5289,16'd2807,-16'd5583,-16'd5496,-16'd6369,-16'd5007,-16'd4859,-16'd1712,16'd2170,-16'd4321,16'd4681};
dout[1105]={ -16'd7843,-16'd674,16'd2990,-16'd2892,-16'd882,16'd3920,-16'd3656,16'd1805,-16'd5778,16'd1522,16'd210,-16'd3956,-16'd7564,16'd4956,16'd4515,-16'd1441,-16'd7635,16'd1853,-16'd4927,-16'd6472,-16'd1918,16'd1879,16'd1467,-16'd4569,16'd7129,-16'd2074,16'd437,-16'd5335,16'd847,-16'd4702,-16'd5468,-16'd3759,-16'd6154,16'd632,-16'd5841,16'd480};
dout[1106]={ 16'd2259,-16'd3132,16'd979,16'd596,-16'd4517,-16'd3136,16'd501,-16'd6039,-16'd5977,-16'd1682,16'd2524,16'd2012,16'd2832,-16'd360,16'd3123,-16'd1833,-16'd6020,16'd2015,-16'd1576,16'd1264,-16'd2067,-16'd4883,16'd4177,16'd3738,-16'd1385,16'd2239,-16'd2964,-16'd4244,-16'd6712,16'd533,16'd2295,-16'd1402,-16'd2695,16'd2289,16'd2899,-16'd9770};
dout[1107]={ 16'd4293,16'd2833,16'd5681,16'd2261,-16'd6378,16'd5779,16'd6047,16'd1323,16'd2058,16'd713,16'd4472,16'd6274,-16'd5556,-16'd6789,16'd3424,16'd4765,-16'd474,-16'd1952,-16'd7252,-16'd2685,16'd4230,-16'd5764,-16'd1957,16'd5600,-16'd675,-16'd775,16'd2825,-16'd188,-16'd1050,16'd6979,16'd7838,16'd2170,16'd1913,16'd2538,16'd1126,-16'd5730};
dout[1108]={ -16'd3447,-16'd490,-16'd263,16'd2207,16'd758,-16'd6082,-16'd6649,16'd8078,16'd2830,16'd2595,-16'd773,16'd5607,16'd793,-16'd3731,16'd6801,16'd4168,-16'd2508,16'd1481,-16'd4235,-16'd4164,16'd5758,-16'd4681,16'd1839,16'd1096,-16'd6187,16'd6185,-16'd5691,-16'd4647,16'd5225,-16'd7821,-16'd2947,16'd3651,-16'd1327,16'd2918,16'd1386,-16'd6559};
dout[1109]={ 16'd1515,16'd1541,16'd6879,-16'd4086,16'd3355,-16'd1576,-16'd1351,16'd3063,16'd7875,16'd2853,16'd3411,-16'd2867,-16'd2608,16'd5574,-16'd5658,-16'd2046,16'd536,16'd1800,16'd2493,16'd2430,16'd3383,16'd3589,-16'd1024,16'd6911,-16'd4960,16'd4950,16'd9208,-16'd5823,16'd4795,16'd6299,-16'd4911,16'd5096,-16'd4068,16'd920,-16'd8441,16'd4828};
dout[1110]={ 16'd775,-16'd3222,-16'd3418,-16'd7583,16'd40,-16'd5160,16'd8537,-16'd10943,-16'd5723,-16'd5649,-16'd2181,-16'd4586,-16'd673,16'd2984,-16'd6902,-16'd2527,16'd5963,16'd3546,-16'd8166,-16'd8630,16'd623,-16'd1917,16'd1216,16'd8379,-16'd13552,16'd452,-16'd1001,16'd7452,-16'd3160,16'd627,16'd6001,-16'd8872,16'd2954,16'd9870,16'd3679,16'd1537};
dout[1111]={ -16'd7508,16'd978,-16'd8468,16'd5308,16'd6690,16'd4271,16'd3100,-16'd6068,-16'd3763,-16'd7329,16'd5686,16'd7535,-16'd2331,-16'd77,-16'd5842,-16'd5395,-16'd3667,-16'd4579,-16'd1022,-16'd2535,-16'd9518,-16'd3861,16'd2160,-16'd7168,-16'd3086,-16'd6181,-16'd2262,16'd1246,16'd424,-16'd6977,16'd3734,16'd1491,-16'd578,16'd1457,-16'd3401,16'd3152};
dout[1112]={ -16'd970,16'd6140,16'd3354,-16'd5643,-16'd2017,16'd5733,16'd5704,-16'd11283,16'd1747,-16'd8819,-16'd8650,-16'd336,-16'd3407,-16'd2417,-16'd6540,-16'd4436,16'd4542,-16'd2039,16'd4406,-16'd4336,-16'd1212,-16'd234,16'd7747,-16'd1129,16'd3809,-16'd7879,16'd2801,-16'd3614,-16'd8168,16'd2993,16'd4901,16'd682,-16'd1302,-16'd7398,16'd2678,-16'd6933};
dout[1113]={ -16'd2243,16'd2084,16'd3853,16'd4557,16'd1272,16'd5616,-16'd4504,-16'd6982,16'd6933,16'd2113,16'd5404,16'd4013,-16'd3511,-16'd5847,-16'd8329,-16'd9464,16'd4592,16'd417,16'd4929,16'd5094,-16'd3414,16'd2894,16'd11,-16'd3178,16'd1854,-16'd4609,16'd2774,16'd3319,-16'd1062,-16'd6980,-16'd1143,-16'd4942,16'd1096,16'd5176,16'd1668,-16'd5854};
dout[1114]={ -16'd7195,-16'd87,16'd7022,16'd974,16'd6996,-16'd8984,16'd2348,-16'd1250,-16'd1733,-16'd7859,16'd6920,-16'd82,-16'd1787,-16'd3675,-16'd7977,16'd2246,16'd2744,-16'd6242,16'd986,-16'd6152,-16'd8291,-16'd9453,-16'd2197,16'd8264,16'd5735,16'd2784,-16'd5424,-16'd2664,16'd2433,-16'd8407,16'd882,-16'd267,-16'd1616,-16'd184,16'd240,-16'd4947};
dout[1115]={ -16'd5408,16'd4302,-16'd5191,16'd2181,-16'd5437,16'd5156,-16'd4203,16'd3032,16'd5429,-16'd3026,-16'd4695,16'd6202,-16'd1660,16'd4378,-16'd8398,-16'd2984,16'd4864,16'd7100,-16'd3658,-16'd4649,16'd4682,-16'd9565,-16'd4137,-16'd3574,16'd1429,-16'd2805,-16'd1945,-16'd8117,16'd1370,16'd3376,16'd1814,-16'd5081,-16'd5973,-16'd5870,16'd142,-16'd7631};
dout[1116]={ 16'd3325,16'd2585,-16'd670,-16'd9387,-16'd235,16'd1731,16'd3833,16'd102,16'd3991,-16'd2519,16'd3578,-16'd804,-16'd3222,16'd3042,-16'd4862,-16'd4021,16'd621,-16'd321,-16'd8508,16'd3096,-16'd959,-16'd5270,-16'd2083,-16'd631,-16'd4356,16'd1587,16'd5601,-16'd2865,-16'd318,16'd2572,-16'd2565,-16'd5299,-16'd2688,16'd4750,-16'd2448,16'd4287};
dout[1117]={ -16'd8585,16'd3889,16'd4074,-16'd3117,-16'd1372,-16'd7722,16'd3764,16'd111,16'd3910,16'd1008,-16'd804,-16'd4563,16'd6194,-16'd5401,16'd909,16'd4350,-16'd1777,16'd2664,16'd994,16'd3010,16'd5011,-16'd4889,-16'd519,-16'd4912,-16'd4386,16'd859,-16'd1287,-16'd3100,-16'd3647,16'd324,-16'd5631,16'd2693,-16'd4094,16'd1391,16'd4517,-16'd2909};
dout[1118]={ -16'd7110,-16'd3760,16'd3208,-16'd618,-16'd2937,-16'd439,16'd7239,-16'd2610,-16'd3906,16'd3959,16'd1104,-16'd480,16'd2353,16'd3462,-16'd4722,-16'd1213,-16'd3613,-16'd824,-16'd4919,-16'd5230,16'd4703,16'd7210,16'd3782,16'd6108,-16'd3438,16'd5895,16'd4111,-16'd613,16'd880,-16'd6762,16'd6946,-16'd2707,-16'd6319,16'd5493,-16'd3392,-16'd4989};
dout[1119]={ -16'd4381,-16'd3543,-16'd3529,-16'd970,-16'd3149,16'd1275,-16'd1581,16'd2864,-16'd1650,16'd4872,16'd3949,16'd2164,16'd4942,16'd5278,-16'd578,-16'd31,-16'd3432,-16'd4208,16'd2716,16'd1269,-16'd6179,16'd2123,-16'd7998,-16'd3556,16'd5412,16'd8315,-16'd4615,-16'd3176,16'd6874,-16'd2013,16'd381,-16'd429,16'd3392,-16'd6759,-16'd505,16'd4628};
dout[1120]={ 16'd1179,16'd785,-16'd1665,-16'd6675,16'd765,-16'd4583,16'd87,-16'd6643,-16'd527,-16'd6578,16'd4838,16'd8771,16'd3167,-16'd1539,16'd6441,-16'd11302,-16'd5067,-16'd5819,-16'd5762,-16'd10375,-16'd6149,16'd2221,-16'd8606,-16'd61,-16'd6880,16'd164,-16'd1453,16'd3949,-16'd7679,-16'd3846,16'd6462,16'd3481,-16'd4150,-16'd2003,-16'd7741,-16'd4911};
dout[1121]={ -16'd7049,-16'd3442,16'd2259,16'd3997,16'd3652,16'd1357,-16'd1835,-16'd2774,16'd2883,-16'd892,16'd2333,-16'd4888,-16'd2488,-16'd7583,16'd939,-16'd4104,-16'd4919,-16'd50,-16'd7992,16'd2250,-16'd5014,16'd5727,-16'd575,-16'd2349,16'd4192,-16'd11145,16'd2331,16'd7912,-16'd7415,-16'd8294,16'd9657,16'd6927,16'd4190,-16'd1492,-16'd2483,-16'd7974};
dout[1122]={ 16'd2871,16'd510,-16'd6842,16'd2729,-16'd3244,16'd5975,-16'd5540,-16'd11100,16'd4001,16'd615,16'd2304,16'd5714,-16'd4823,-16'd9413,16'd635,-16'd6029,-16'd7267,-16'd2941,-16'd5967,-16'd8750,-16'd4266,-16'd2624,-16'd6319,16'd5575,16'd3427,-16'd9744,16'd5528,-16'd363,-16'd6507,-16'd5266,16'd7762,16'd7092,-16'd8750,-16'd10788,-16'd318,16'd6832};
dout[1123]={ -16'd8320,-16'd646,-16'd4816,-16'd1337,16'd551,-16'd6805,-16'd6920,-16'd5020,-16'd2239,-16'd7068,-16'd5488,16'd1491,16'd9185,-16'd4731,-16'd1018,-16'd739,16'd4492,16'd3281,-16'd8236,-16'd31,16'd1521,16'd1005,16'd4141,-16'd377,-16'd704,-16'd7493,-16'd8182,16'd6353,-16'd2219,16'd2425,-16'd11157,16'd3690,16'd2394,-16'd810,16'd1328,-16'd5672};
dout[1124]={ -16'd5770,16'd1189,-16'd3493,-16'd4772,-16'd2054,-16'd7410,-16'd2291,-16'd4394,16'd1323,-16'd9367,-16'd5647,16'd3147,16'd1670,16'd6835,-16'd5561,16'd1211,16'd4077,16'd225,-16'd6245,-16'd3144,-16'd8160,-16'd1366,-16'd688,16'd7941,16'd2196,-16'd7049,-16'd7192,16'd3506,16'd4715,16'd6576,-16'd7305,-16'd3549,-16'd2436,16'd3948,-16'd3567,-16'd5337};
dout[1125]={ -16'd9267,16'd3494,16'd617,-16'd7315,16'd4400,16'd5143,16'd2104,-16'd7632,16'd2457,-16'd718,16'd4815,-16'd3756,16'd4770,16'd1029,16'd1557,-16'd1833,16'd1001,-16'd3772,-16'd2125,16'd2134,16'd5608,-16'd2881,16'd3639,16'd2307,16'd5706,16'd2116,16'd7421,16'd989,-16'd7027,-16'd7988,-16'd6564,16'd4455,-16'd2606,16'd5837,-16'd6035,16'd7173};
dout[1126]={ 16'd1598,16'd22,16'd6029,-16'd8013,16'd2645,16'd5350,-16'd2487,16'd6371,16'd4640,-16'd796,-16'd5384,16'd8013,-16'd294,-16'd3689,-16'd6114,16'd7984,-16'd4392,-16'd168,16'd3373,16'd2198,-16'd6193,-16'd2835,-16'd4568,-16'd648,-16'd3630,-16'd1044,-16'd5485,-16'd1969,-16'd272,16'd2962,-16'd3741,16'd3282,-16'd7740,-16'd95,16'd4658,-16'd6242};
dout[1127]={ 16'd4997,-16'd1393,16'd5730,16'd6976,16'd1359,-16'd7022,16'd481,-16'd112,-16'd9143,16'd2735,-16'd576,-16'd3578,-16'd6369,16'd2696,-16'd46,16'd4421,-16'd5360,-16'd1809,16'd4006,16'd2035,16'd2238,16'd1234,16'd4355,-16'd1947,16'd5079,16'd3175,16'd289,16'd675,-16'd5820,-16'd3352,16'd5413,16'd3236,-16'd6329,-16'd5935,-16'd8194,-16'd4955};
dout[1128]={ -16'd6065,16'd2931,-16'd2159,-16'd4236,-16'd1131,16'd5982,-16'd805,-16'd3675,-16'd737,-16'd1476,-16'd2548,16'd1811,16'd4245,-16'd3772,-16'd2765,16'd3916,-16'd7720,-16'd205,-16'd3256,-16'd2253,16'd1975,-16'd4086,-16'd6470,-16'd4088,-16'd8609,16'd7834,16'd6695,-16'd4626,-16'd2705,-16'd2719,-16'd5597,-16'd2616,16'd5478,-16'd4035,-16'd2269,-16'd5968};
dout[1129]={ -16'd2391,16'd3962,-16'd102,-16'd3714,16'd3013,16'd2534,16'd6418,16'd10316,-16'd7036,-16'd3481,-16'd5647,-16'd138,16'd6831,-16'd1254,16'd3884,16'd7169,-16'd619,16'd4654,16'd5388,-16'd1811,-16'd1651,16'd8533,-16'd4840,-16'd73,16'd528,-16'd3166,-16'd3126,-16'd7161,-16'd3237,16'd241,16'd5061,16'd2840,-16'd777,16'd2868,16'd662,16'd4257};
dout[1130]={ 16'd2105,16'd1223,-16'd1618,-16'd8246,16'd2306,-16'd1963,16'd5966,-16'd11518,-16'd10195,16'd3072,16'd4255,16'd7393,-16'd2330,-16'd4560,16'd5889,-16'd33,-16'd9003,16'd2350,16'd1097,16'd2379,-16'd3726,16'd4489,-16'd4036,16'd925,-16'd4428,-16'd10132,16'd8503,16'd7589,-16'd3407,16'd179,16'd2847,-16'd1790,-16'd4355,-16'd3267,-16'd2589,16'd4242};
dout[1131]={ 16'd2201,16'd3219,-16'd9681,-16'd3132,16'd6913,16'd6087,-16'd5766,-16'd5076,-16'd7159,-16'd6653,-16'd6656,16'd5334,16'd8370,16'd5557,16'd215,-16'd1456,16'd1068,-16'd9131,16'd2021,16'd4360,16'd1096,16'd4717,-16'd2725,16'd5634,-16'd6093,-16'd6506,-16'd6797,-16'd4623,-16'd4649,-16'd5114,16'd2866,16'd4359,-16'd5214,-16'd4558,-16'd2069,-16'd7193};
dout[1132]={ 16'd6505,16'd8638,-16'd9555,16'd3365,-16'd4118,-16'd4895,-16'd1462,16'd4273,16'd1584,-16'd6060,-16'd7056,-16'd4885,-16'd4003,16'd3611,16'd7770,-16'd1295,16'd185,-16'd788,16'd313,-16'd6753,-16'd10127,-16'd5894,16'd4823,16'd2568,16'd380,-16'd10465,16'd3468,16'd2122,-16'd8677,-16'd6738,16'd7417,-16'd3199,-16'd8684,-16'd13178,16'd612,16'd4480};
dout[1133]={ 16'd4096,16'd1264,16'd6072,-16'd4174,-16'd1755,-16'd4120,16'd583,-16'd5681,16'd8955,-16'd5471,-16'd3704,16'd6435,16'd8412,16'd4999,16'd85,-16'd2785,-16'd4443,16'd5087,-16'd9679,16'd4356,-16'd1805,-16'd5828,-16'd5300,16'd5793,16'd11249,16'd2307,16'd2721,16'd6430,16'd3517,-16'd7581,-16'd6460,-16'd102,-16'd2174,-16'd7611,-16'd1749,16'd3176};
dout[1134]={ 16'd523,16'd4618,-16'd5887,16'd2919,-16'd649,-16'd4053,-16'd623,16'd4763,-16'd5641,-16'd10173,16'd6420,-16'd1951,16'd6957,-16'd5517,-16'd6631,-16'd28,-16'd6537,-16'd5422,16'd2770,-16'd4696,16'd2265,16'd2949,-16'd5491,16'd1148,-16'd4499,-16'd1991,-16'd2816,-16'd5159,-16'd1459,-16'd4696,-16'd7955,16'd3143,-16'd7756,16'd6423,-16'd1213,-16'd2589};
dout[1135]={ -16'd4342,-16'd7300,16'd3624,16'd3909,-16'd1928,-16'd6816,-16'd5511,-16'd7779,16'd5444,16'd3855,16'd1299,-16'd2129,16'd2574,-16'd2529,16'd3819,16'd1185,16'd5369,16'd704,-16'd1948,-16'd6915,16'd6770,-16'd5746,16'd4510,16'd2593,16'd6799,16'd4827,-16'd1710,-16'd3389,-16'd2186,-16'd65,16'd3711,16'd3827,-16'd482,16'd3785,-16'd3262,16'd394};
dout[1136]={ -16'd9076,16'd151,-16'd3539,16'd3779,-16'd2967,-16'd7597,-16'd1975,-16'd6264,-16'd3800,-16'd6609,-16'd3886,16'd1960,16'd8309,-16'd2576,-16'd2702,16'd341,-16'd1585,16'd6436,-16'd3240,-16'd3144,-16'd6140,-16'd8065,-16'd8074,-16'd3723,-16'd301,-16'd1576,16'd5679,16'd5910,-16'd7549,-16'd3621,16'd2698,16'd4634,-16'd6527,16'd3934,-16'd9280,16'd2203};
dout[1137]={ 16'd4662,16'd4368,-16'd5503,-16'd1137,16'd804,16'd4504,-16'd3224,16'd1943,16'd18,16'd160,-16'd6679,-16'd4922,16'd7430,-16'd675,16'd5948,16'd283,-16'd6617,-16'd4763,-16'd5510,16'd3409,16'd2482,16'd1990,-16'd4566,16'd2958,-16'd1029,16'd5042,-16'd8370,-16'd1701,-16'd979,-16'd3871,16'd2665,-16'd4748,-16'd4020,-16'd1657,-16'd106,-16'd5889};
dout[1138]={ -16'd1742,-16'd1698,-16'd3427,16'd3678,16'd3729,16'd7428,16'd1690,16'd4819,16'd5006,16'd1348,-16'd5729,16'd681,16'd2857,16'd7795,-16'd7738,16'd5414,-16'd6516,16'd3073,-16'd8347,16'd4046,16'd4689,16'd2099,16'd3684,16'd6590,16'd3526,16'd794,16'd4239,16'd945,16'd4523,-16'd3071,-16'd4857,-16'd8011,16'd92,-16'd5233,16'd1060,-16'd4958};
dout[1139]={ 16'd6685,-16'd4397,16'd1782,16'd1927,-16'd4553,16'd145,-16'd1177,-16'd894,16'd2475,16'd6367,-16'd4686,-16'd5734,-16'd1750,16'd712,-16'd6690,-16'd3254,16'd1823,-16'd3645,16'd2321,16'd2792,16'd1454,16'd4712,16'd1500,16'd859,-16'd6349,16'd1764,-16'd9402,-16'd3589,-16'd746,-16'd1964,-16'd1166,16'd4119,16'd1972,16'd6204,16'd3596,16'd3322};
dout[1140]={ -16'd4298,16'd4995,-16'd6741,16'd2510,16'd9303,-16'd4105,-16'd1693,-16'd137,-16'd1265,16'd565,16'd9831,-16'd1741,16'd7761,-16'd9904,16'd2512,-16'd6297,-16'd6855,-16'd4674,-16'd3144,-16'd8271,16'd28,-16'd8442,16'd40,16'd6619,-16'd5592,-16'd2918,16'd5560,16'd1283,-16'd1970,16'd4167,16'd1977,16'd7312,-16'd6897,-16'd11898,-16'd3754,16'd5791};
dout[1141]={ 16'd3024,-16'd2693,16'd587,-16'd5955,16'd1853,16'd4909,16'd3776,-16'd3964,-16'd4106,-16'd5460,-16'd8270,16'd4442,-16'd1437,-16'd3958,16'd425,16'd5739,-16'd5020,-16'd8325,-16'd969,-16'd7225,-16'd2399,-16'd6290,16'd863,-16'd3770,16'd1190,16'd275,16'd5853,16'd4861,-16'd10008,16'd2124,16'd367,-16'd6350,-16'd2878,-16'd7364,16'd3489,-16'd2226};
dout[1142]={ -16'd7269,-16'd4568,-16'd8769,-16'd4650,-16'd3883,16'd4003,16'd3638,-16'd2629,16'd4510,16'd2259,-16'd9572,-16'd3290,-16'd4718,-16'd3797,-16'd4498,16'd224,-16'd5282,-16'd7505,16'd3539,16'd6590,-16'd2131,-16'd7092,-16'd218,16'd2203,16'd6724,16'd1109,16'd2529,16'd1074,-16'd3126,-16'd9659,16'd3313,16'd312,-16'd4454,-16'd6823,16'd6344,-16'd5112};
dout[1143]={ -16'd2742,-16'd126,16'd5020,-16'd6038,16'd5802,-16'd5580,-16'd7409,16'd2288,-16'd656,16'd3986,-16'd1362,-16'd5166,-16'd3307,-16'd6547,-16'd4887,16'd7803,16'd3177,16'd622,16'd2053,16'd6208,-16'd7190,-16'd9884,-16'd7565,16'd3003,16'd3419,-16'd10114,16'd2602,16'd4737,16'd5632,-16'd5286,-16'd12385,16'd4563,-16'd4075,-16'd3244,-16'd2011,-16'd4538};
dout[1144]={ 16'd7050,16'd5240,-16'd410,-16'd7779,16'd1914,-16'd5476,16'd4479,16'd821,-16'd2058,16'd2249,16'd5305,16'd3989,-16'd2302,16'd171,16'd4395,16'd2580,-16'd6653,-16'd1430,-16'd1912,-16'd2431,-16'd4968,-16'd8258,-16'd1672,-16'd4545,-16'd1194,16'd4102,-16'd2210,16'd4847,-16'd774,-16'd2426,-16'd5566,16'd1042,16'd4036,-16'd7344,-16'd328,16'd2781};
dout[1145]={ -16'd189,-16'd6342,16'd6663,16'd5122,16'd3083,-16'd1069,16'd718,-16'd9402,16'd1338,-16'd2749,16'd7323,16'd239,16'd3855,16'd1781,16'd4016,-16'd3946,-16'd4305,16'd7295,-16'd5877,16'd5975,-16'd2322,-16'd4362,-16'd1402,16'd538,-16'd825,-16'd2698,16'd5914,16'd2416,-16'd2423,16'd6817,-16'd2712,16'd2328,-16'd1582,16'd940,16'd3945,-16'd162};
dout[1146]={ 16'd4859,16'd286,16'd3558,16'd3163,-16'd2346,-16'd5275,-16'd1955,16'd2210,16'd870,16'd3470,-16'd5595,-16'd2667,16'd439,16'd3096,-16'd7650,16'd5778,-16'd6972,-16'd1484,-16'd5862,-16'd7497,16'd5413,-16'd677,16'd160,16'd2753,16'd895,16'd2186,-16'd5829,-16'd377,-16'd6079,16'd3137,-16'd1557,-16'd703,16'd5812,16'd1700,-16'd6152,-16'd2334};
dout[1147]={ -16'd2744,-16'd4161,-16'd5767,16'd3129,16'd2450,-16'd5699,16'd5256,16'd2999,16'd1533,-16'd4585,16'd3000,16'd4311,16'd3343,-16'd5247,-16'd1865,-16'd2687,-16'd4189,-16'd5575,16'd3533,16'd1575,-16'd5358,16'd2278,16'd4890,-16'd5851,16'd1077,-16'd303,-16'd7153,16'd3527,16'd1714,16'd946,-16'd4520,16'd1762,-16'd2530,-16'd181,-16'd1590,-16'd7032};
dout[1148]={ -16'd3668,16'd1061,16'd5456,16'd699,16'd5195,-16'd2847,16'd1632,16'd7189,16'd2580,16'd4996,16'd7014,-16'd3021,16'd4186,-16'd883,-16'd1011,16'd6907,-16'd6513,-16'd6597,16'd7046,-16'd7842,-16'd7883,16'd2686,16'd6394,-16'd4700,-16'd731,-16'd5356,16'd1106,-16'd5031,16'd5555,16'd10878,-16'd5,16'd4304,16'd1665,-16'd3613,16'd2452,-16'd4515};
dout[1149]={ -16'd5411,16'd4962,16'd3946,16'd4050,-16'd3834,16'd2757,16'd4956,-16'd299,-16'd1426,16'd4414,-16'd4533,16'd3886,-16'd5396,-16'd5215,-16'd3720,-16'd6614,16'd4122,16'd3136,-16'd2863,16'd6021,-16'd3094,-16'd2939,16'd5619,-16'd920,-16'd7341,16'd8011,-16'd7731,-16'd9520,16'd2087,-16'd198,16'd1201,16'd953,-16'd4346,16'd847,-16'd7133,16'd5970};
dout[1150]={ -16'd4929,-16'd8102,16'd4107,16'd2943,-16'd3138,-16'd2639,-16'd133,16'd1969,16'd282,16'd6095,16'd582,-16'd4151,16'd779,-16'd9373,16'd3079,-16'd8548,-16'd1310,16'd7346,-16'd1275,-16'd103,16'd4548,-16'd3831,16'd98,16'd7306,-16'd1855,16'd1607,16'd3016,16'd5317,-16'd8005,16'd911,16'd4292,-16'd6487,-16'd6143,-16'd9508,16'd3881,16'd4728};
dout[1151]={ 16'd1858,16'd215,-16'd5154,16'd665,-16'd5053,16'd8328,-16'd5900,-16'd2625,-16'd1543,16'd5220,16'd5389,-16'd2624,16'd347,-16'd2950,16'd1571,-16'd5087,-16'd1234,-16'd5744,-16'd3517,16'd5897,-16'd522,16'd1628,16'd4745,-16'd4019,-16'd8824,-16'd1372,-16'd4681,16'd5902,-16'd5254,16'd3012,16'd12113,-16'd5202,-16'd2562,-16'd8933,16'd8741,-16'd8206};
dout[1152]={ -16'd2136,16'd5014,-16'd6496,-16'd5194,16'd2043,-16'd4070,16'd2847,16'd7147,-16'd1519,16'd4195,-16'd7637,-16'd2514,16'd754,16'd387,-16'd4862,16'd1327,-16'd4850,-16'd6560,-16'd3342,-16'd6097,16'd2676,-16'd9902,16'd8398,16'd4200,16'd4262,-16'd3678,16'd7271,-16'd7533,-16'd4385,16'd5407,16'd3085,-16'd8038,16'd5186,-16'd3217,-16'd1890,16'd3267};
dout[1153]={ -16'd617,-16'd3282,16'd3435,16'd2534,16'd6712,16'd35,-16'd3173,16'd4165,16'd7830,16'd3970,16'd6146,16'd4107,-16'd3992,16'd3388,16'd622,-16'd3713,-16'd1867,-16'd3925,-16'd4482,16'd493,16'd4437,-16'd7591,16'd3053,16'd3870,-16'd2639,-16'd4903,-16'd3227,16'd4293,-16'd7653,16'd5344,-16'd12404,-16'd6202,16'd1595,-16'd8979,-16'd4276,-16'd1220};
dout[1154]={ -16'd4388,16'd3991,-16'd4740,16'd5184,16'd7974,-16'd4550,-16'd1725,16'd3603,-16'd1379,-16'd5945,-16'd1592,16'd1089,16'd3978,-16'd6119,-16'd1327,-16'd4393,-16'd4027,16'd3126,-16'd540,16'd4013,-16'd402,-16'd8860,-16'd6690,16'd7369,-16'd2529,-16'd5989,16'd3835,-16'd5787,-16'd4781,16'd3665,-16'd5520,-16'd1774,16'd911,-16'd3636,-16'd4546,16'd3875};
dout[1155]={ -16'd4423,-16'd1907,16'd1047,-16'd3192,16'd5855,-16'd2297,16'd6002,16'd1782,-16'd3378,-16'd6667,16'd966,-16'd1001,16'd6829,16'd156,16'd4988,16'd6384,16'd7499,-16'd1682,16'd7392,16'd2233,16'd7725,-16'd6483,-16'd6344,-16'd1044,-16'd433,-16'd3400,16'd7842,-16'd2981,-16'd4790,-16'd5910,-16'd6885,-16'd7742,16'd514,16'd5676,16'd5426,-16'd5597};
dout[1156]={ 16'd2852,-16'd4036,-16'd976,-16'd3993,16'd2623,16'd1106,16'd1854,-16'd2077,-16'd5920,-16'd5821,16'd867,16'd734,-16'd3725,-16'd3635,-16'd1006,16'd7629,-16'd370,-16'd3540,-16'd5241,16'd3306,-16'd1188,-16'd5926,-16'd4410,16'd1390,-16'd4429,16'd295,-16'd4673,-16'd5298,-16'd3563,-16'd6217,-16'd913,-16'd4215,-16'd2889,-16'd1475,16'd585,-16'd6322};
dout[1157]={ 16'd1389,-16'd5943,-16'd5779,-16'd48,16'd4135,16'd534,-16'd7255,-16'd4968,-16'd685,16'd3771,-16'd7741,-16'd2507,16'd3244,16'd1123,16'd5731,16'd1471,-16'd7542,16'd6629,-16'd3721,16'd4570,16'd1705,16'd7028,-16'd3422,16'd6350,-16'd9499,-16'd442,-16'd3687,-16'd6583,16'd1265,16'd6778,-16'd1657,16'd3042,16'd7398,-16'd3795,-16'd5096,16'd3244};
dout[1158]={ 16'd2717,16'd3206,16'd6185,-16'd1666,16'd5035,-16'd6584,-16'd6058,-16'd4803,16'd510,16'd3360,16'd4273,-16'd342,-16'd4384,-16'd1185,-16'd684,16'd5224,-16'd4191,16'd2173,16'd433,-16'd1768,16'd3179,16'd265,-16'd268,-16'd5606,-16'd3069,16'd5755,-16'd7036,-16'd7526,-16'd8311,-16'd547,16'd6835,-16'd2205,16'd5130,-16'd5176,16'd4894,16'd6786};
dout[1159]={ 16'd4249,16'd2148,-16'd5504,16'd7477,-16'd5167,-16'd6781,-16'd5940,16'd6232,16'd7428,-16'd256,16'd1741,16'd6723,-16'd2279,16'd1928,-16'd4541,-16'd3052,16'd4405,-16'd2997,-16'd5636,-16'd5910,-16'd4008,16'd5419,-16'd1943,-16'd1345,-16'd7433,16'd6402,-16'd7390,-16'd4034,-16'd8182,16'd9947,16'd1743,16'd99,16'd6977,-16'd2660,-16'd6466,16'd3345};
dout[1160]={ -16'd3721,-16'd116,-16'd7995,-16'd2674,16'd2085,-16'd398,-16'd7828,16'd6810,16'd903,-16'd2666,16'd4801,-16'd94,16'd4337,-16'd9321,-16'd3258,16'd6820,-16'd3827,16'd9224,-16'd6927,-16'd8865,-16'd4987,-16'd5142,-16'd2992,16'd771,-16'd1017,-16'd7227,16'd8323,-16'd7987,16'd1985,16'd2427,16'd8730,-16'd3783,-16'd5740,-16'd3400,16'd1809,-16'd6127};
dout[1161]={ 16'd2007,-16'd10303,16'd5122,16'd1391,16'd7264,16'd1514,-16'd5098,16'd4595,16'd5646,16'd3425,-16'd6843,-16'd2005,16'd3931,-16'd2066,16'd7114,16'd5942,-16'd5488,-16'd2750,-16'd9276,-16'd4057,-16'd1641,-16'd7826,16'd8002,-16'd80,-16'd10364,-16'd3251,-16'd2596,-16'd3078,16'd3506,-16'd8212,-16'd2327,-16'd5388,-16'd6733,16'd3671,-16'd3751,16'd5414};
dout[1162]={ -16'd8520,-16'd4010,-16'd1062,-16'd4497,-16'd9050,-16'd8197,-16'd1029,16'd1111,16'd3093,16'd3204,-16'd4410,16'd1577,-16'd1673,16'd2625,16'd2217,16'd2453,16'd5777,16'd6838,16'd617,16'd2284,16'd6382,16'd441,-16'd4352,16'd7023,-16'd2028,16'd2393,16'd2,-16'd3014,16'd445,16'd297,-16'd2391,16'd552,16'd1153,-16'd4487,16'd4342,16'd4516};
dout[1163]={ 16'd5615,-16'd3383,16'd7495,16'd1919,-16'd5901,-16'd949,-16'd4912,-16'd5511,16'd7347,16'd8120,16'd6905,16'd112,-16'd2732,-16'd1421,16'd3115,16'd2691,-16'd8529,16'd620,-16'd886,-16'd4542,16'd5197,-16'd8050,16'd3695,-16'd7523,16'd2159,-16'd160,16'd655,16'd376,-16'd3668,-16'd5093,-16'd1969,16'd2568,16'd1963,16'd5328,16'd4683,-16'd6913};
dout[1164]={ -16'd7271,-16'd6336,16'd3239,-16'd5143,16'd8016,16'd2399,16'd1782,-16'd6830,-16'd4216,16'd3458,16'd66,16'd3492,16'd6302,16'd4549,16'd1229,16'd1806,-16'd1430,16'd7201,-16'd1775,16'd7425,16'd4972,-16'd5901,16'd6282,-16'd7646,-16'd1734,16'd2875,-16'd1828,16'd2594,16'd1401,-16'd3305,-16'd10673,-16'd3035,16'd4524,16'd259,-16'd2929,-16'd2088};
dout[1165]={ -16'd3222,16'd1848,-16'd5540,-16'd4608,-16'd3253,-16'd4452,-16'd2614,16'd1834,16'd2696,-16'd6223,16'd4523,16'd1371,16'd2966,16'd5310,16'd4855,-16'd611,16'd1178,-16'd1742,-16'd2222,16'd7071,-16'd2722,-16'd1432,-16'd2497,16'd5753,-16'd3202,-16'd80,-16'd4491,-16'd1115,16'd5431,16'd5786,16'd6953,-16'd5431,16'd4127,-16'd2566,-16'd2874,-16'd2069};
dout[1166]={ 16'd5010,16'd1963,-16'd4588,16'd6248,16'd2472,16'd958,-16'd7555,-16'd3351,16'd6062,-16'd6561,16'd4920,-16'd3744,-16'd6558,-16'd2035,16'd189,-16'd2622,16'd510,16'd1567,16'd2904,-16'd225,16'd2178,-16'd831,-16'd5827,-16'd4099,-16'd4480,-16'd3557,-16'd4931,-16'd2914,-16'd6904,-16'd2132,-16'd1614,-16'd3831,16'd3670,16'd6415,16'd2418,-16'd6514};
dout[1167]={ 16'd1933,-16'd5341,-16'd6284,-16'd2581,-16'd3621,16'd293,-16'd7302,-16'd7918,16'd6822,16'd599,-16'd2352,-16'd6858,16'd5515,16'd8109,-16'd4688,16'd868,-16'd5603,-16'd3242,16'd5043,-16'd2695,16'd172,-16'd3802,-16'd3908,16'd1686,16'd1875,16'd7501,16'd5630,-16'd7606,-16'd9563,16'd5586,16'd2350,16'd1410,16'd7245,-16'd2825,16'd5365,16'd5911};
dout[1168]={ 16'd6052,-16'd522,16'd4327,16'd6686,16'd4514,-16'd4177,16'd3578,-16'd3595,16'd4732,-16'd3494,16'd4178,16'd183,16'd4255,-16'd2429,-16'd8171,-16'd2960,16'd3080,16'd5961,16'd501,16'd4198,-16'd1922,16'd1706,-16'd4636,-16'd6354,-16'd4842,16'd2396,-16'd5355,-16'd6673,16'd1448,16'd706,16'd422,-16'd1624,-16'd7451,16'd8760,-16'd2740,-16'd892};
dout[1169]={ -16'd7053,16'd6218,16'd3424,-16'd2186,-16'd3926,-16'd1984,-16'd3799,-16'd558,16'd4078,-16'd824,16'd5576,16'd1810,16'd2628,-16'd4810,-16'd3612,16'd668,-16'd3826,-16'd4713,16'd1516,-16'd723,-16'd7076,-16'd4118,-16'd2151,-16'd1093,16'd2732,16'd4193,-16'd8300,-16'd7264,16'd182,-16'd4795,-16'd1910,16'd5415,-16'd5699,-16'd988,16'd5059,16'd9590};
dout[1170]={ 16'd1119,16'd502,16'd5443,16'd2776,16'd32,-16'd1769,16'd425,16'd1151,16'd707,16'd4758,-16'd373,-16'd5581,16'd9817,16'd4913,-16'd4589,-16'd800,-16'd5778,16'd3705,-16'd6354,-16'd8037,16'd784,-16'd5710,-16'd2834,16'd7655,-16'd9441,-16'd2068,16'd7638,-16'd8666,16'd3723,16'd4529,16'd221,-16'd4291,-16'd242,-16'd11813,16'd8366,-16'd6788};
dout[1171]={ 16'd3639,-16'd10002,-16'd598,-16'd6936,-16'd212,-16'd1017,16'd5474,-16'd6666,16'd7120,-16'd6325,16'd2617,16'd7326,-16'd6988,-16'd6710,16'd4088,-16'd2090,16'd5883,-16'd472,-16'd5051,-16'd7673,16'd1316,-16'd9054,16'd7036,16'd4024,16'd1203,-16'd3732,-16'd2831,16'd5310,16'd5264,-16'd4722,16'd8693,16'd1917,-16'd6322,-16'd1775,16'd5091,16'd3153};
dout[1172]={ -16'd7350,16'd4744,-16'd4772,-16'd302,16'd2179,-16'd5511,16'd3974,16'd8041,16'd7756,16'd1320,-16'd5283,16'd3145,-16'd5412,-16'd2486,16'd3494,16'd2299,16'd4610,16'd5380,16'd268,16'd5679,16'd653,16'd2981,16'd8010,-16'd6967,-16'd7844,-16'd6915,16'd6807,16'd3819,16'd460,-16'd8776,16'd5417,16'd1333,-16'd4523,-16'd1138,-16'd6754,-16'd3493};
dout[1173]={ 16'd4050,-16'd4110,-16'd4116,16'd8335,16'd2783,16'd4209,16'd1923,16'd8411,-16'd5239,16'd161,-16'd1788,16'd3068,-16'd1046,-16'd2952,16'd3393,-16'd7485,16'd254,16'd6219,-16'd8340,-16'd1216,16'd2335,-16'd10768,16'd17,-16'd3679,16'd3452,-16'd6752,-16'd2870,-16'd6957,-16'd2402,-16'd4784,-16'd11781,-16'd2014,-16'd1989,-16'd739,16'd5876,16'd1389};
dout[1174]={ -16'd1793,16'd3867,16'd6560,-16'd1442,16'd1309,-16'd6771,16'd343,16'd3524,-16'd699,16'd126,-16'd4269,16'd5230,-16'd852,-16'd3895,-16'd5831,16'd155,-16'd248,16'd6362,-16'd5314,16'd915,-16'd4308,-16'd939,-16'd6467,-16'd8146,16'd1666,16'd6113,-16'd4150,-16'd319,-16'd6683,-16'd7766,-16'd8781,-16'd4438,16'd6344,16'd3221,-16'd6268,16'd6158};
dout[1175]={ -16'd1854,16'd6456,-16'd6441,-16'd1406,-16'd2277,-16'd3655,16'd61,-16'd6735,-16'd1767,16'd2835,16'd1505,-16'd4130,-16'd4038,16'd5840,-16'd2033,-16'd6623,16'd910,16'd1250,16'd5966,-16'd3991,-16'd5781,-16'd7136,-16'd7338,16'd5581,16'd3190,-16'd6757,-16'd5058,16'd2847,-16'd5334,-16'd7310,-16'd6331,16'd3145,16'd2815,16'd4180,-16'd5645,16'd469};
dout[1176]={ -16'd666,16'd4235,16'd3455,-16'd5705,16'd7982,-16'd3556,16'd1379,16'd4176,-16'd4297,16'd4661,-16'd2657,16'd1457,16'd3150,-16'd7227,-16'd8286,-16'd1673,16'd479,16'd1794,16'd4002,-16'd2523,-16'd1838,-16'd6059,16'd4674,16'd5398,16'd1474,-16'd2464,16'd4831,-16'd2786,-16'd2387,16'd2347,16'd5959,-16'd7107,16'd850,-16'd2578,16'd1980,16'd5289};
dout[1177]={ -16'd2950,-16'd3501,-16'd2820,16'd1714,16'd2235,-16'd102,16'd7325,-16'd1119,16'd324,16'd392,-16'd4157,16'd4189,-16'd2308,16'd6805,16'd5426,16'd2731,16'd747,16'd5307,16'd4631,-16'd48,16'd5236,16'd1462,-16'd4443,16'd1310,-16'd2556,16'd3293,-16'd3310,-16'd176,16'd3451,-16'd5589,-16'd3655,16'd1904,-16'd6203,16'd218,-16'd6199,-16'd2570};
dout[1178]={ 16'd4807,16'd7625,-16'd1498,16'd2733,16'd82,-16'd7679,-16'd5063,-16'd4056,-16'd5635,-16'd5331,-16'd2311,16'd4775,-16'd4285,-16'd1839,-16'd1246,16'd1622,-16'd6389,16'd351,-16'd3366,-16'd6015,-16'd113,16'd6221,-16'd65,-16'd6215,-16'd4607,16'd1482,-16'd3479,-16'd1362,-16'd7109,16'd6349,-16'd1822,-16'd4988,-16'd5282,-16'd2682,-16'd981,-16'd5460};
dout[1179]={ -16'd8311,-16'd3434,-16'd2675,16'd1998,16'd4401,16'd547,16'd5540,16'd2339,-16'd1041,16'd5491,16'd6195,-16'd5664,-16'd4189,-16'd1032,16'd7148,16'd3607,-16'd6018,-16'd3070,16'd626,-16'd644,16'd1345,-16'd1159,16'd4577,16'd3470,-16'd1613,16'd6214,-16'd11554,16'd2300,16'd4326,16'd1595,16'd3300,16'd4022,16'd6548,16'd142,16'd4368,-16'd3384};
dout[1180]={ -16'd4264,16'd817,16'd3778,-16'd7247,-16'd3680,16'd2907,-16'd9377,16'd1057,-16'd7449,-16'd7385,16'd5492,-16'd1956,16'd2889,-16'd3555,-16'd3780,16'd1199,16'd2948,16'd2483,-16'd6175,16'd3755,-16'd1949,-16'd9061,16'd5336,16'd6797,-16'd45,-16'd1186,-16'd4542,-16'd6741,16'd3415,-16'd2888,-16'd248,-16'd5649,16'd7152,-16'd7948,-16'd1131,-16'd6537};
dout[1181]={ -16'd514,-16'd7148,16'd6664,16'd7096,-16'd7554,-16'd5179,16'd5171,16'd6555,16'd1563,-16'd1317,-16'd4931,16'd3596,16'd9396,16'd1576,16'd4771,-16'd4101,-16'd3339,16'd4107,16'd4467,-16'd5168,-16'd3952,-16'd148,16'd4104,-16'd5574,16'd1671,-16'd6273,-16'd3504,16'd802,-16'd6361,16'd1120,-16'd4013,16'd4893,-16'd3332,16'd2836,16'd858,16'd3489};
dout[1182]={ -16'd1307,-16'd1737,-16'd5835,16'd1689,16'd1603,16'd213,-16'd4246,16'd3006,-16'd3109,16'd3835,16'd5169,-16'd537,16'd4883,16'd3766,16'd2718,-16'd2808,16'd5070,16'd4884,16'd2949,-16'd3650,-16'd4899,-16'd3960,16'd5844,-16'd8481,-16'd8474,-16'd7418,-16'd2639,-16'd2597,-16'd4736,16'd845,-16'd4726,-16'd1553,16'd955,16'd6759,16'd132,16'd4193};
dout[1183]={ -16'd6689,-16'd2707,-16'd8850,-16'd1415,16'd2952,16'd3859,16'd564,-16'd3376,-16'd6254,16'd2651,16'd3809,-16'd6403,-16'd6109,16'd4493,-16'd6494,-16'd7134,-16'd2749,16'd7118,-16'd4020,-16'd4475,16'd1769,-16'd1630,-16'd2214,-16'd11181,16'd4836,-16'd689,-16'd1526,-16'd8318,-16'd5922,16'd2665,-16'd5224,16'd2317,-16'd2927,-16'd1607,16'd1106,16'd5364};
dout[1184]={ -16'd6597,16'd6973,16'd5522,-16'd1404,-16'd5754,16'd5651,16'd963,16'd1503,-16'd1285,16'd8170,-16'd5449,16'd4311,16'd4475,16'd517,-16'd6337,16'd4518,16'd865,-16'd4199,16'd2582,-16'd6235,16'd3081,-16'd39,16'd6023,16'd2443,16'd5094,16'd2013,16'd3603,16'd438,-16'd1495,16'd1588,-16'd2287,-16'd6500,-16'd3349,-16'd2688,-16'd3696,16'd3714};
dout[1185]={ -16'd353,16'd707,16'd2994,-16'd1824,16'd4818,16'd3380,-16'd2821,-16'd1249,-16'd3094,-16'd3142,16'd282,-16'd5784,-16'd588,-16'd4090,16'd6608,16'd382,-16'd992,16'd3988,-16'd7370,-16'd636,-16'd5613,16'd338,-16'd702,-16'd7659,-16'd2476,-16'd7425,-16'd1641,-16'd6240,16'd6539,16'd4413,16'd5959,16'd824,16'd4910,-16'd412,16'd3728,-16'd2768};
dout[1186]={ 16'd4569,-16'd5237,-16'd2442,-16'd5294,-16'd1970,16'd456,-16'd4976,16'd6166,16'd1500,16'd3349,-16'd2549,-16'd3939,-16'd5284,16'd6253,-16'd8154,-16'd4047,16'd6055,-16'd3759,-16'd390,-16'd4806,16'd3741,16'd481,16'd7855,-16'd5768,16'd978,-16'd7184,16'd4370,-16'd8719,-16'd518,16'd2811,16'd1552,-16'd7163,16'd4890,16'd6574,16'd233,16'd4599};
dout[1187]={ -16'd1844,16'd4152,16'd4909,-16'd567,16'd3363,-16'd2823,-16'd5429,-16'd1515,16'd4485,16'd635,-16'd7623,16'd606,16'd3607,-16'd618,-16'd3224,-16'd238,-16'd4703,16'd7290,-16'd709,16'd6265,16'd7125,16'd5316,-16'd3753,-16'd4882,-16'd4427,-16'd4187,-16'd8969,-16'd6768,-16'd2699,-16'd4137,-16'd1229,16'd1809,-16'd6499,16'd6349,16'd1918,16'd2606};
dout[1188]={ -16'd5763,-16'd622,16'd1596,-16'd2080,16'd5703,16'd6458,16'd707,16'd2018,16'd885,16'd285,-16'd1472,-16'd3093,16'd1494,16'd7486,16'd633,-16'd1666,16'd4721,-16'd2848,16'd54,16'd6571,16'd96,16'd3301,-16'd5927,-16'd3721,16'd5146,-16'd4414,16'd1888,16'd2843,-16'd6147,16'd3227,16'd519,16'd5685,-16'd104,16'd539,16'd161,16'd4721};
dout[1189]={ 16'd1955,16'd4575,16'd2769,16'd2625,-16'd5753,16'd6078,-16'd4939,16'd2920,-16'd1148,-16'd1597,16'd6519,16'd8460,16'd3280,16'd4123,16'd4695,16'd5148,-16'd855,-16'd4360,16'd3637,-16'd5227,16'd2921,16'd3454,-16'd4775,16'd6964,-16'd2053,-16'd1897,-16'd12977,-16'd2238,16'd4377,16'd2126,16'd2350,16'd1914,-16'd7201,16'd321,-16'd3763,16'd4441};
dout[1190]={ 16'd4217,16'd2988,-16'd4415,-16'd2817,-16'd1192,16'd4020,-16'd1352,16'd8211,16'd760,-16'd7317,-16'd5523,16'd2181,16'd5993,-16'd1881,16'd2534,-16'd3821,16'd2844,16'd6135,-16'd6010,16'd4232,16'd466,-16'd5482,16'd2427,16'd8033,16'd3735,16'd7145,16'd726,16'd3216,-16'd1298,16'd2174,16'd9895,-16'd8548,16'd2867,16'd521,-16'd865,-16'd128};
dout[1191]={ -16'd4630,16'd4022,-16'd8449,-16'd8776,16'd2301,16'd298,16'd2766,16'd3033,-16'd4401,16'd2923,-16'd1222,16'd1701,16'd2407,-16'd7305,-16'd1174,16'd6538,16'd3614,-16'd2826,16'd2872,-16'd1608,-16'd2216,-16'd122,-16'd5630,16'd1205,-16'd764,-16'd5915,16'd1098,16'd3728,-16'd594,-16'd7431,-16'd4188,-16'd619,-16'd4903,16'd5315,16'd6606,-16'd2593};
dout[1192]={ -16'd5580,16'd2694,-16'd7492,16'd2055,-16'd3716,16'd6313,-16'd4792,16'd7300,16'd3084,16'd2803,-16'd1969,16'd5284,16'd3821,16'd611,-16'd1548,16'd193,-16'd2044,-16'd8043,-16'd3269,16'd2180,-16'd4650,16'd2336,16'd2273,16'd3435,-16'd456,-16'd1470,16'd249,16'd356,-16'd7981,-16'd9797,16'd1274,16'd2978,-16'd1070,16'd4759,16'd4424,-16'd3246};
dout[1193]={ 16'd4047,-16'd3176,-16'd3328,-16'd6824,-16'd1594,16'd5264,16'd4313,16'd4696,16'd3209,-16'd2193,16'd2868,16'd7023,-16'd3170,16'd992,-16'd3875,16'd5951,-16'd5802,16'd2473,-16'd1124,-16'd2902,-16'd2745,16'd351,-16'd3787,-16'd2739,-16'd4142,-16'd3367,16'd2013,-16'd1197,16'd193,16'd2429,-16'd6018,16'd6788,16'd3721,-16'd6029,16'd1718,16'd1596};
dout[1194]={ -16'd2438,16'd6,16'd2593,16'd4207,-16'd347,16'd6639,16'd2201,16'd872,16'd2032,16'd4896,-16'd2002,16'd5597,16'd1158,-16'd7435,-16'd2302,-16'd8170,16'd1700,-16'd4875,-16'd3342,-16'd6013,-16'd6963,16'd3610,16'd5263,-16'd11247,-16'd5383,16'd1173,-16'd1554,-16'd6713,-16'd4331,-16'd3955,16'd341,16'd3126,16'd5318,16'd3011,-16'd1331,16'd1207};
dout[1195]={ 16'd5445,16'd1837,-16'd7291,16'd1552,16'd8340,16'd5982,16'd1087,-16'd987,16'd605,16'd1074,16'd729,-16'd2171,-16'd1941,16'd6596,-16'd6396,16'd5265,-16'd8168,16'd7311,16'd804,-16'd4879,16'd1690,16'd3473,16'd4571,16'd4038,16'd7477,-16'd3993,16'd3346,16'd201,16'd6010,-16'd7686,-16'd5437,-16'd1706,-16'd3385,16'd5914,-16'd9779,-16'd1747};
dout[1196]={ 16'd5033,16'd2779,-16'd5984,16'd1883,16'd5401,-16'd4438,-16'd4393,16'd2590,-16'd480,-16'd2718,16'd1277,16'd4911,-16'd3891,16'd2107,16'd1619,16'd1035,16'd1921,16'd3660,-16'd4025,16'd5339,-16'd5078,-16'd722,16'd3437,16'd5247,-16'd3168,16'd6637,-16'd6036,16'd1530,16'd5499,16'd1745,16'd1109,16'd5113,-16'd3782,-16'd2965,-16'd1507,16'd5445};
dout[1197]={ -16'd789,16'd1438,16'd4342,-16'd2150,-16'd3629,16'd1317,16'd7019,-16'd5296,-16'd4034,-16'd795,16'd7032,16'd3863,16'd8229,16'd1465,-16'd2719,16'd5046,-16'd46,16'd1270,16'd6572,16'd5618,16'd2645,-16'd5967,16'd5008,16'd3580,-16'd4841,16'd5186,16'd1031,-16'd3403,16'd1937,16'd2915,16'd2471,16'd2397,-16'd8013,16'd1870,-16'd8042,16'd3154};
dout[1198]={ 16'd3347,-16'd303,16'd3967,-16'd2317,16'd1340,-16'd3548,-16'd365,-16'd3766,-16'd985,16'd9170,16'd22,-16'd2702,-16'd166,-16'd4875,-16'd1970,16'd1238,16'd4132,-16'd4128,16'd4521,-16'd343,-16'd5672,-16'd6507,-16'd4420,16'd4095,-16'd4249,-16'd3345,-16'd7026,-16'd3369,-16'd6309,16'd1753,-16'd3302,16'd3442,16'd3049,16'd3065,16'd2285,-16'd2589};
dout[1199]={ -16'd1388,16'd2971,16'd1426,-16'd5810,16'd3441,-16'd3358,16'd2597,16'd1195,-16'd5292,-16'd468,-16'd164,16'd6362,16'd9738,16'd4154,16'd3251,-16'd7370,16'd4785,-16'd4311,16'd7888,16'd768,16'd5396,-16'd2002,16'd8695,-16'd5784,-16'd4948,16'd6140,16'd863,16'd4206,-16'd4604,16'd5527,-16'd2852,-16'd7711,16'd6131,16'd458,-16'd6593,-16'd467};
end     
always @ (posedge clk) begin

w <= dout[addr];
end

endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */
